
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e8",x"de",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e8",x"de",x"c2"),
    14 => (x"48",x"e8",x"cc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c6",x"dc"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"48",x"72",x"4c"),
    72 => (x"7c",x"70",x"98",x"ff"),
    73 => (x"bf",x"e8",x"cc",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"ff",x"c3",x"48",x"71"),
    79 => (x"d0",x"7c",x"70",x"98"),
    80 => (x"29",x"d0",x"49",x"66"),
    81 => (x"ff",x"c3",x"48",x"71"),
    82 => (x"d0",x"7c",x"70",x"98"),
    83 => (x"29",x"c8",x"49",x"66"),
    84 => (x"ff",x"c3",x"48",x"71"),
    85 => (x"d0",x"7c",x"70",x"98"),
    86 => (x"ff",x"c3",x"48",x"66"),
    87 => (x"72",x"7c",x"70",x"98"),
    88 => (x"71",x"29",x"d0",x"49"),
    89 => (x"98",x"ff",x"c3",x"48"),
    90 => (x"4b",x"6c",x"7c",x"70"),
    91 => (x"4d",x"ff",x"f0",x"c9"),
    92 => (x"05",x"ab",x"ff",x"c3"),
    93 => (x"ff",x"c3",x"87",x"d0"),
    94 => (x"c1",x"4b",x"6c",x"7c"),
    95 => (x"87",x"c6",x"02",x"8d"),
    96 => (x"02",x"ab",x"ff",x"c3"),
    97 => (x"48",x"73",x"87",x"f0"),
    98 => (x"1e",x"87",x"ff",x"fd"),
    99 => (x"d4",x"ff",x"49",x"c0"),
   100 => (x"78",x"ff",x"c3",x"48"),
   101 => (x"c8",x"c3",x"81",x"c1"),
   102 => (x"f1",x"04",x"a9",x"b7"),
   103 => (x"1e",x"4f",x"26",x"87"),
   104 => (x"87",x"e7",x"1e",x"73"),
   105 => (x"4b",x"df",x"f8",x"c4"),
   106 => (x"ff",x"c0",x"1e",x"c0"),
   107 => (x"49",x"f7",x"c1",x"f0"),
   108 => (x"c4",x"87",x"df",x"fd"),
   109 => (x"05",x"a8",x"c1",x"86"),
   110 => (x"ff",x"87",x"ea",x"c0"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c0",x"c0",x"c1",x"78"),
   113 => (x"1e",x"c0",x"c0",x"c0"),
   114 => (x"c1",x"f0",x"e1",x"c0"),
   115 => (x"c1",x"fd",x"49",x"e9"),
   116 => (x"70",x"86",x"c4",x"87"),
   117 => (x"87",x"ca",x"05",x"98"),
   118 => (x"c3",x"48",x"d4",x"ff"),
   119 => (x"48",x"c1",x"78",x"ff"),
   120 => (x"e6",x"fe",x"87",x"cb"),
   121 => (x"05",x"8b",x"c1",x"87"),
   122 => (x"c0",x"87",x"fd",x"fe"),
   123 => (x"87",x"de",x"fc",x"48"),
   124 => (x"ff",x"1e",x"73",x"1e"),
   125 => (x"ff",x"c3",x"48",x"d4"),
   126 => (x"c0",x"4b",x"d3",x"78"),
   127 => (x"f0",x"ff",x"c0",x"1e"),
   128 => (x"fc",x"49",x"c1",x"c1"),
   129 => (x"86",x"c4",x"87",x"cc"),
   130 => (x"ca",x"05",x"98",x"70"),
   131 => (x"48",x"d4",x"ff",x"87"),
   132 => (x"c1",x"78",x"ff",x"c3"),
   133 => (x"fd",x"87",x"cb",x"48"),
   134 => (x"8b",x"c1",x"87",x"f1"),
   135 => (x"87",x"db",x"ff",x"05"),
   136 => (x"e9",x"fb",x"48",x"c0"),
   137 => (x"5b",x"5e",x"0e",x"87"),
   138 => (x"d4",x"ff",x"0e",x"5c"),
   139 => (x"87",x"db",x"fd",x"4c"),
   140 => (x"c0",x"1e",x"ea",x"c6"),
   141 => (x"c8",x"c1",x"f0",x"e1"),
   142 => (x"87",x"d6",x"fb",x"49"),
   143 => (x"a8",x"c1",x"86",x"c4"),
   144 => (x"fe",x"87",x"c8",x"02"),
   145 => (x"48",x"c0",x"87",x"ea"),
   146 => (x"fa",x"87",x"e2",x"c1"),
   147 => (x"49",x"70",x"87",x"d2"),
   148 => (x"99",x"ff",x"ff",x"cf"),
   149 => (x"02",x"a9",x"ea",x"c6"),
   150 => (x"d3",x"fe",x"87",x"c8"),
   151 => (x"c1",x"48",x"c0",x"87"),
   152 => (x"ff",x"c3",x"87",x"cb"),
   153 => (x"4b",x"f1",x"c0",x"7c"),
   154 => (x"70",x"87",x"f4",x"fc"),
   155 => (x"eb",x"c0",x"02",x"98"),
   156 => (x"c0",x"1e",x"c0",x"87"),
   157 => (x"fa",x"c1",x"f0",x"ff"),
   158 => (x"87",x"d6",x"fa",x"49"),
   159 => (x"98",x"70",x"86",x"c4"),
   160 => (x"c3",x"87",x"d9",x"05"),
   161 => (x"49",x"6c",x"7c",x"ff"),
   162 => (x"7c",x"7c",x"ff",x"c3"),
   163 => (x"c0",x"c1",x"7c",x"7c"),
   164 => (x"87",x"c4",x"02",x"99"),
   165 => (x"87",x"d5",x"48",x"c1"),
   166 => (x"87",x"d1",x"48",x"c0"),
   167 => (x"c4",x"05",x"ab",x"c2"),
   168 => (x"c8",x"48",x"c0",x"87"),
   169 => (x"05",x"8b",x"c1",x"87"),
   170 => (x"c0",x"87",x"fd",x"fe"),
   171 => (x"87",x"dc",x"f9",x"48"),
   172 => (x"c2",x"1e",x"73",x"1e"),
   173 => (x"c1",x"48",x"e8",x"cc"),
   174 => (x"ff",x"4b",x"c7",x"78"),
   175 => (x"78",x"c2",x"48",x"d0"),
   176 => (x"ff",x"87",x"c8",x"fb"),
   177 => (x"78",x"c3",x"48",x"d0"),
   178 => (x"e5",x"c0",x"1e",x"c0"),
   179 => (x"49",x"c0",x"c1",x"d0"),
   180 => (x"c4",x"87",x"ff",x"f8"),
   181 => (x"05",x"a8",x"c1",x"86"),
   182 => (x"c2",x"4b",x"87",x"c1"),
   183 => (x"87",x"c5",x"05",x"ab"),
   184 => (x"f9",x"c0",x"48",x"c0"),
   185 => (x"05",x"8b",x"c1",x"87"),
   186 => (x"fc",x"87",x"d0",x"ff"),
   187 => (x"cc",x"c2",x"87",x"f7"),
   188 => (x"98",x"70",x"58",x"ec"),
   189 => (x"c1",x"87",x"cd",x"05"),
   190 => (x"f0",x"ff",x"c0",x"1e"),
   191 => (x"f8",x"49",x"d0",x"c1"),
   192 => (x"86",x"c4",x"87",x"d0"),
   193 => (x"c3",x"48",x"d4",x"ff"),
   194 => (x"fd",x"c2",x"78",x"ff"),
   195 => (x"f0",x"cc",x"c2",x"87"),
   196 => (x"48",x"d0",x"ff",x"58"),
   197 => (x"d4",x"ff",x"78",x"c2"),
   198 => (x"78",x"ff",x"c3",x"48"),
   199 => (x"ed",x"f7",x"48",x"c1"),
   200 => (x"5b",x"5e",x"0e",x"87"),
   201 => (x"71",x"0e",x"5d",x"5c"),
   202 => (x"c5",x"4c",x"c0",x"4b"),
   203 => (x"4a",x"df",x"cd",x"ee"),
   204 => (x"c3",x"48",x"d4",x"ff"),
   205 => (x"48",x"68",x"78",x"ff"),
   206 => (x"05",x"a8",x"fe",x"c3"),
   207 => (x"ff",x"87",x"fe",x"c0"),
   208 => (x"9b",x"73",x"4d",x"d4"),
   209 => (x"d0",x"87",x"cc",x"02"),
   210 => (x"49",x"73",x"1e",x"66"),
   211 => (x"c4",x"87",x"e8",x"f5"),
   212 => (x"ff",x"87",x"d6",x"86"),
   213 => (x"d1",x"c4",x"48",x"d0"),
   214 => (x"7d",x"ff",x"c3",x"78"),
   215 => (x"c1",x"48",x"66",x"d0"),
   216 => (x"58",x"a6",x"d4",x"88"),
   217 => (x"f0",x"05",x"98",x"70"),
   218 => (x"48",x"d4",x"ff",x"87"),
   219 => (x"78",x"78",x"ff",x"c3"),
   220 => (x"c5",x"05",x"9b",x"73"),
   221 => (x"48",x"d0",x"ff",x"87"),
   222 => (x"4a",x"c1",x"78",x"d0"),
   223 => (x"05",x"8a",x"c1",x"4c"),
   224 => (x"74",x"87",x"ed",x"fe"),
   225 => (x"87",x"c2",x"f6",x"48"),
   226 => (x"71",x"1e",x"73",x"1e"),
   227 => (x"ff",x"4b",x"c0",x"4a"),
   228 => (x"ff",x"c3",x"48",x"d4"),
   229 => (x"48",x"d0",x"ff",x"78"),
   230 => (x"ff",x"78",x"c3",x"c4"),
   231 => (x"ff",x"c3",x"48",x"d4"),
   232 => (x"c0",x"1e",x"72",x"78"),
   233 => (x"d1",x"c1",x"f0",x"ff"),
   234 => (x"87",x"e6",x"f5",x"49"),
   235 => (x"98",x"70",x"86",x"c4"),
   236 => (x"c8",x"87",x"d2",x"05"),
   237 => (x"66",x"cc",x"1e",x"c0"),
   238 => (x"87",x"e5",x"fd",x"49"),
   239 => (x"4b",x"70",x"86",x"c4"),
   240 => (x"c2",x"48",x"d0",x"ff"),
   241 => (x"f5",x"48",x"73",x"78"),
   242 => (x"5e",x"0e",x"87",x"c4"),
   243 => (x"0e",x"5d",x"5c",x"5b"),
   244 => (x"ff",x"c0",x"1e",x"c0"),
   245 => (x"49",x"c9",x"c1",x"f0"),
   246 => (x"d2",x"87",x"f7",x"f4"),
   247 => (x"f0",x"cc",x"c2",x"1e"),
   248 => (x"87",x"fd",x"fc",x"49"),
   249 => (x"4c",x"c0",x"86",x"c8"),
   250 => (x"b7",x"d2",x"84",x"c1"),
   251 => (x"87",x"f8",x"04",x"ac"),
   252 => (x"97",x"f0",x"cc",x"c2"),
   253 => (x"c0",x"c3",x"49",x"bf"),
   254 => (x"a9",x"c0",x"c1",x"99"),
   255 => (x"87",x"e7",x"c0",x"05"),
   256 => (x"97",x"f7",x"cc",x"c2"),
   257 => (x"31",x"d0",x"49",x"bf"),
   258 => (x"97",x"f8",x"cc",x"c2"),
   259 => (x"32",x"c8",x"4a",x"bf"),
   260 => (x"cc",x"c2",x"b1",x"72"),
   261 => (x"4a",x"bf",x"97",x"f9"),
   262 => (x"cf",x"4c",x"71",x"b1"),
   263 => (x"9c",x"ff",x"ff",x"ff"),
   264 => (x"34",x"ca",x"84",x"c1"),
   265 => (x"c2",x"87",x"e7",x"c1"),
   266 => (x"bf",x"97",x"f9",x"cc"),
   267 => (x"c6",x"31",x"c1",x"49"),
   268 => (x"fa",x"cc",x"c2",x"99"),
   269 => (x"c7",x"4a",x"bf",x"97"),
   270 => (x"b1",x"72",x"2a",x"b7"),
   271 => (x"97",x"f5",x"cc",x"c2"),
   272 => (x"cf",x"4d",x"4a",x"bf"),
   273 => (x"f6",x"cc",x"c2",x"9d"),
   274 => (x"c3",x"4a",x"bf",x"97"),
   275 => (x"c2",x"32",x"ca",x"9a"),
   276 => (x"bf",x"97",x"f7",x"cc"),
   277 => (x"73",x"33",x"c2",x"4b"),
   278 => (x"f8",x"cc",x"c2",x"b2"),
   279 => (x"c3",x"4b",x"bf",x"97"),
   280 => (x"b7",x"c6",x"9b",x"c0"),
   281 => (x"c2",x"b2",x"73",x"2b"),
   282 => (x"71",x"48",x"c1",x"81"),
   283 => (x"c1",x"49",x"70",x"30"),
   284 => (x"70",x"30",x"75",x"48"),
   285 => (x"c1",x"4c",x"72",x"4d"),
   286 => (x"c8",x"94",x"71",x"84"),
   287 => (x"06",x"ad",x"b7",x"c0"),
   288 => (x"34",x"c1",x"87",x"cc"),
   289 => (x"c0",x"c8",x"2d",x"b7"),
   290 => (x"ff",x"01",x"ad",x"b7"),
   291 => (x"48",x"74",x"87",x"f4"),
   292 => (x"0e",x"87",x"f7",x"f1"),
   293 => (x"5d",x"5c",x"5b",x"5e"),
   294 => (x"c2",x"86",x"f8",x"0e"),
   295 => (x"c0",x"48",x"d6",x"d5"),
   296 => (x"ce",x"cd",x"c2",x"78"),
   297 => (x"fb",x"49",x"c0",x"1e"),
   298 => (x"86",x"c4",x"87",x"de"),
   299 => (x"c5",x"05",x"98",x"70"),
   300 => (x"c9",x"48",x"c0",x"87"),
   301 => (x"4d",x"c0",x"87",x"c0"),
   302 => (x"ed",x"c0",x"7e",x"c1"),
   303 => (x"c2",x"49",x"bf",x"e6"),
   304 => (x"71",x"4a",x"c4",x"ce"),
   305 => (x"e0",x"ee",x"4b",x"c8"),
   306 => (x"05",x"98",x"70",x"87"),
   307 => (x"7e",x"c0",x"87",x"c2"),
   308 => (x"bf",x"e2",x"ed",x"c0"),
   309 => (x"e0",x"ce",x"c2",x"49"),
   310 => (x"4b",x"c8",x"71",x"4a"),
   311 => (x"70",x"87",x"ca",x"ee"),
   312 => (x"87",x"c2",x"05",x"98"),
   313 => (x"02",x"6e",x"7e",x"c0"),
   314 => (x"c2",x"87",x"fd",x"c0"),
   315 => (x"4d",x"bf",x"d4",x"d4"),
   316 => (x"9f",x"cc",x"d5",x"c2"),
   317 => (x"c5",x"48",x"7e",x"bf"),
   318 => (x"05",x"a8",x"ea",x"d6"),
   319 => (x"d4",x"c2",x"87",x"c7"),
   320 => (x"ce",x"4d",x"bf",x"d4"),
   321 => (x"ca",x"48",x"6e",x"87"),
   322 => (x"02",x"a8",x"d5",x"e9"),
   323 => (x"48",x"c0",x"87",x"c5"),
   324 => (x"c2",x"87",x"e3",x"c7"),
   325 => (x"75",x"1e",x"ce",x"cd"),
   326 => (x"87",x"ec",x"f9",x"49"),
   327 => (x"98",x"70",x"86",x"c4"),
   328 => (x"c0",x"87",x"c5",x"05"),
   329 => (x"87",x"ce",x"c7",x"48"),
   330 => (x"bf",x"e2",x"ed",x"c0"),
   331 => (x"e0",x"ce",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f2",x"ec"),
   334 => (x"87",x"c8",x"05",x"98"),
   335 => (x"48",x"d6",x"d5",x"c2"),
   336 => (x"87",x"da",x"78",x"c1"),
   337 => (x"bf",x"e6",x"ed",x"c0"),
   338 => (x"c4",x"ce",x"c2",x"49"),
   339 => (x"4b",x"c8",x"71",x"4a"),
   340 => (x"70",x"87",x"d6",x"ec"),
   341 => (x"c5",x"c0",x"02",x"98"),
   342 => (x"c6",x"48",x"c0",x"87"),
   343 => (x"d5",x"c2",x"87",x"d8"),
   344 => (x"49",x"bf",x"97",x"cc"),
   345 => (x"05",x"a9",x"d5",x"c1"),
   346 => (x"c2",x"87",x"cd",x"c0"),
   347 => (x"bf",x"97",x"cd",x"d5"),
   348 => (x"a9",x"ea",x"c2",x"49"),
   349 => (x"87",x"c5",x"c0",x"02"),
   350 => (x"f9",x"c5",x"48",x"c0"),
   351 => (x"ce",x"cd",x"c2",x"87"),
   352 => (x"48",x"7e",x"bf",x"97"),
   353 => (x"02",x"a8",x"e9",x"c3"),
   354 => (x"6e",x"87",x"ce",x"c0"),
   355 => (x"a8",x"eb",x"c3",x"48"),
   356 => (x"87",x"c5",x"c0",x"02"),
   357 => (x"dd",x"c5",x"48",x"c0"),
   358 => (x"d9",x"cd",x"c2",x"87"),
   359 => (x"99",x"49",x"bf",x"97"),
   360 => (x"87",x"cc",x"c0",x"05"),
   361 => (x"97",x"da",x"cd",x"c2"),
   362 => (x"a9",x"c2",x"49",x"bf"),
   363 => (x"87",x"c5",x"c0",x"02"),
   364 => (x"c1",x"c5",x"48",x"c0"),
   365 => (x"db",x"cd",x"c2",x"87"),
   366 => (x"c2",x"48",x"bf",x"97"),
   367 => (x"70",x"58",x"d2",x"d5"),
   368 => (x"88",x"c1",x"48",x"4c"),
   369 => (x"58",x"d6",x"d5",x"c2"),
   370 => (x"97",x"dc",x"cd",x"c2"),
   371 => (x"81",x"75",x"49",x"bf"),
   372 => (x"97",x"dd",x"cd",x"c2"),
   373 => (x"32",x"c8",x"4a",x"bf"),
   374 => (x"c2",x"7e",x"a1",x"72"),
   375 => (x"6e",x"48",x"e3",x"d9"),
   376 => (x"de",x"cd",x"c2",x"78"),
   377 => (x"c8",x"48",x"bf",x"97"),
   378 => (x"d5",x"c2",x"58",x"a6"),
   379 => (x"c2",x"02",x"bf",x"d6"),
   380 => (x"ed",x"c0",x"87",x"cf"),
   381 => (x"c2",x"49",x"bf",x"e2"),
   382 => (x"71",x"4a",x"e0",x"ce"),
   383 => (x"e8",x"e9",x"4b",x"c8"),
   384 => (x"02",x"98",x"70",x"87"),
   385 => (x"c0",x"87",x"c5",x"c0"),
   386 => (x"87",x"ea",x"c3",x"48"),
   387 => (x"bf",x"ce",x"d5",x"c2"),
   388 => (x"f7",x"d9",x"c2",x"4c"),
   389 => (x"f3",x"cd",x"c2",x"5c"),
   390 => (x"c8",x"49",x"bf",x"97"),
   391 => (x"f2",x"cd",x"c2",x"31"),
   392 => (x"a1",x"4a",x"bf",x"97"),
   393 => (x"f4",x"cd",x"c2",x"49"),
   394 => (x"d0",x"4a",x"bf",x"97"),
   395 => (x"49",x"a1",x"72",x"32"),
   396 => (x"97",x"f5",x"cd",x"c2"),
   397 => (x"32",x"d8",x"4a",x"bf"),
   398 => (x"c4",x"49",x"a1",x"72"),
   399 => (x"d9",x"c2",x"91",x"66"),
   400 => (x"c2",x"81",x"bf",x"e3"),
   401 => (x"c2",x"59",x"eb",x"d9"),
   402 => (x"bf",x"97",x"fb",x"cd"),
   403 => (x"c2",x"32",x"c8",x"4a"),
   404 => (x"bf",x"97",x"fa",x"cd"),
   405 => (x"c2",x"4a",x"a2",x"4b"),
   406 => (x"bf",x"97",x"fc",x"cd"),
   407 => (x"73",x"33",x"d0",x"4b"),
   408 => (x"cd",x"c2",x"4a",x"a2"),
   409 => (x"4b",x"bf",x"97",x"fd"),
   410 => (x"33",x"d8",x"9b",x"cf"),
   411 => (x"c2",x"4a",x"a2",x"73"),
   412 => (x"c2",x"5a",x"ef",x"d9"),
   413 => (x"c2",x"92",x"74",x"8a"),
   414 => (x"72",x"48",x"ef",x"d9"),
   415 => (x"c1",x"c1",x"78",x"a1"),
   416 => (x"e0",x"cd",x"c2",x"87"),
   417 => (x"c8",x"49",x"bf",x"97"),
   418 => (x"df",x"cd",x"c2",x"31"),
   419 => (x"a1",x"4a",x"bf",x"97"),
   420 => (x"c7",x"31",x"c5",x"49"),
   421 => (x"29",x"c9",x"81",x"ff"),
   422 => (x"59",x"f7",x"d9",x"c2"),
   423 => (x"97",x"e5",x"cd",x"c2"),
   424 => (x"32",x"c8",x"4a",x"bf"),
   425 => (x"97",x"e4",x"cd",x"c2"),
   426 => (x"4a",x"a2",x"4b",x"bf"),
   427 => (x"6e",x"92",x"66",x"c4"),
   428 => (x"f3",x"d9",x"c2",x"82"),
   429 => (x"eb",x"d9",x"c2",x"5a"),
   430 => (x"c2",x"78",x"c0",x"48"),
   431 => (x"72",x"48",x"e7",x"d9"),
   432 => (x"d9",x"c2",x"78",x"a1"),
   433 => (x"d9",x"c2",x"48",x"f7"),
   434 => (x"c2",x"78",x"bf",x"eb"),
   435 => (x"c2",x"48",x"fb",x"d9"),
   436 => (x"78",x"bf",x"ef",x"d9"),
   437 => (x"bf",x"d6",x"d5",x"c2"),
   438 => (x"87",x"c9",x"c0",x"02"),
   439 => (x"30",x"c4",x"48",x"74"),
   440 => (x"c9",x"c0",x"7e",x"70"),
   441 => (x"f3",x"d9",x"c2",x"87"),
   442 => (x"30",x"c4",x"48",x"bf"),
   443 => (x"d5",x"c2",x"7e",x"70"),
   444 => (x"78",x"6e",x"48",x"da"),
   445 => (x"8e",x"f8",x"48",x"c1"),
   446 => (x"4c",x"26",x"4d",x"26"),
   447 => (x"4f",x"26",x"4b",x"26"),
   448 => (x"5c",x"5b",x"5e",x"0e"),
   449 => (x"4a",x"71",x"0e",x"5d"),
   450 => (x"bf",x"d6",x"d5",x"c2"),
   451 => (x"72",x"87",x"cb",x"02"),
   452 => (x"72",x"2b",x"c7",x"4b"),
   453 => (x"9d",x"ff",x"c1",x"4d"),
   454 => (x"4b",x"72",x"87",x"c9"),
   455 => (x"4d",x"72",x"2b",x"c8"),
   456 => (x"c2",x"9d",x"ff",x"c3"),
   457 => (x"83",x"bf",x"e3",x"d9"),
   458 => (x"bf",x"de",x"ed",x"c0"),
   459 => (x"87",x"d9",x"02",x"ab"),
   460 => (x"5b",x"e2",x"ed",x"c0"),
   461 => (x"1e",x"ce",x"cd",x"c2"),
   462 => (x"cb",x"f1",x"49",x"73"),
   463 => (x"70",x"86",x"c4",x"87"),
   464 => (x"87",x"c5",x"05",x"98"),
   465 => (x"e6",x"c0",x"48",x"c0"),
   466 => (x"d6",x"d5",x"c2",x"87"),
   467 => (x"87",x"d2",x"02",x"bf"),
   468 => (x"91",x"c4",x"49",x"75"),
   469 => (x"81",x"ce",x"cd",x"c2"),
   470 => (x"ff",x"cf",x"4c",x"69"),
   471 => (x"9c",x"ff",x"ff",x"ff"),
   472 => (x"49",x"75",x"87",x"cb"),
   473 => (x"cd",x"c2",x"91",x"c2"),
   474 => (x"69",x"9f",x"81",x"ce"),
   475 => (x"fe",x"48",x"74",x"4c"),
   476 => (x"5e",x"0e",x"87",x"c6"),
   477 => (x"0e",x"5d",x"5c",x"5b"),
   478 => (x"4c",x"71",x"86",x"f8"),
   479 => (x"87",x"c5",x"05",x"9c"),
   480 => (x"c0",x"c3",x"48",x"c0"),
   481 => (x"7e",x"a4",x"c8",x"87"),
   482 => (x"d8",x"78",x"c0",x"48"),
   483 => (x"87",x"c7",x"02",x"66"),
   484 => (x"bf",x"97",x"66",x"d8"),
   485 => (x"c0",x"87",x"c5",x"05"),
   486 => (x"87",x"e9",x"c2",x"48"),
   487 => (x"49",x"c1",x"1e",x"c0"),
   488 => (x"87",x"e3",x"c7",x"49"),
   489 => (x"4d",x"70",x"86",x"c4"),
   490 => (x"c2",x"c1",x"02",x"9d"),
   491 => (x"de",x"d5",x"c2",x"87"),
   492 => (x"49",x"66",x"d8",x"4a"),
   493 => (x"70",x"87",x"d7",x"e2"),
   494 => (x"f2",x"c0",x"02",x"98"),
   495 => (x"d8",x"4a",x"75",x"87"),
   496 => (x"4b",x"cb",x"49",x"66"),
   497 => (x"70",x"87",x"fc",x"e2"),
   498 => (x"e2",x"c0",x"02",x"98"),
   499 => (x"75",x"1e",x"c0",x"87"),
   500 => (x"87",x"c7",x"02",x"9d"),
   501 => (x"c0",x"48",x"a6",x"c8"),
   502 => (x"c8",x"87",x"c5",x"78"),
   503 => (x"78",x"c1",x"48",x"a6"),
   504 => (x"c6",x"49",x"66",x"c8"),
   505 => (x"86",x"c4",x"87",x"e1"),
   506 => (x"05",x"9d",x"4d",x"70"),
   507 => (x"75",x"87",x"fe",x"fe"),
   508 => (x"ce",x"c1",x"02",x"9d"),
   509 => (x"49",x"a5",x"dc",x"87"),
   510 => (x"78",x"69",x"48",x"6e"),
   511 => (x"c4",x"49",x"a5",x"da"),
   512 => (x"a4",x"c4",x"48",x"a6"),
   513 => (x"48",x"69",x"9f",x"78"),
   514 => (x"78",x"08",x"66",x"c4"),
   515 => (x"bf",x"d6",x"d5",x"c2"),
   516 => (x"d4",x"87",x"d2",x"02"),
   517 => (x"69",x"9f",x"49",x"a5"),
   518 => (x"ff",x"ff",x"c0",x"49"),
   519 => (x"d0",x"48",x"71",x"99"),
   520 => (x"c2",x"7e",x"70",x"30"),
   521 => (x"6e",x"7e",x"c0",x"87"),
   522 => (x"bf",x"66",x"c4",x"48"),
   523 => (x"08",x"66",x"c4",x"80"),
   524 => (x"cc",x"7c",x"c0",x"78"),
   525 => (x"66",x"c4",x"49",x"a4"),
   526 => (x"a4",x"d0",x"79",x"bf"),
   527 => (x"c1",x"79",x"c0",x"49"),
   528 => (x"c0",x"87",x"c2",x"48"),
   529 => (x"fa",x"8e",x"f8",x"48"),
   530 => (x"5e",x"0e",x"87",x"ee"),
   531 => (x"71",x"0e",x"5c",x"5b"),
   532 => (x"c1",x"02",x"9c",x"4c"),
   533 => (x"a4",x"c8",x"87",x"cb"),
   534 => (x"c1",x"02",x"69",x"49"),
   535 => (x"49",x"6c",x"87",x"c3"),
   536 => (x"71",x"48",x"66",x"cc"),
   537 => (x"58",x"a6",x"d0",x"80"),
   538 => (x"d5",x"c2",x"b9",x"70"),
   539 => (x"ff",x"4a",x"bf",x"d2"),
   540 => (x"71",x"99",x"72",x"ba"),
   541 => (x"e5",x"c0",x"02",x"99"),
   542 => (x"4b",x"a4",x"c4",x"87"),
   543 => (x"ff",x"f9",x"49",x"6b"),
   544 => (x"c2",x"7b",x"70",x"87"),
   545 => (x"49",x"bf",x"ce",x"d5"),
   546 => (x"7c",x"71",x"81",x"6c"),
   547 => (x"c2",x"b9",x"66",x"cc"),
   548 => (x"4a",x"bf",x"d2",x"d5"),
   549 => (x"99",x"72",x"ba",x"ff"),
   550 => (x"ff",x"05",x"99",x"71"),
   551 => (x"66",x"cc",x"87",x"db"),
   552 => (x"87",x"d6",x"f9",x"7c"),
   553 => (x"71",x"1e",x"73",x"1e"),
   554 => (x"c7",x"02",x"9b",x"4b"),
   555 => (x"49",x"a3",x"c8",x"87"),
   556 => (x"87",x"c5",x"05",x"69"),
   557 => (x"f6",x"c0",x"48",x"c0"),
   558 => (x"e7",x"d9",x"c2",x"87"),
   559 => (x"a3",x"c4",x"49",x"bf"),
   560 => (x"c2",x"4a",x"6a",x"4a"),
   561 => (x"ce",x"d5",x"c2",x"8a"),
   562 => (x"a1",x"72",x"92",x"bf"),
   563 => (x"d2",x"d5",x"c2",x"49"),
   564 => (x"9a",x"6b",x"4a",x"bf"),
   565 => (x"c0",x"49",x"a1",x"72"),
   566 => (x"c8",x"59",x"e2",x"ed"),
   567 => (x"ea",x"71",x"1e",x"66"),
   568 => (x"86",x"c4",x"87",x"e6"),
   569 => (x"c4",x"05",x"98",x"70"),
   570 => (x"c2",x"48",x"c0",x"87"),
   571 => (x"f8",x"48",x"c1",x"87"),
   572 => (x"73",x"1e",x"87",x"ca"),
   573 => (x"9b",x"4b",x"71",x"1e"),
   574 => (x"87",x"e4",x"c0",x"02"),
   575 => (x"5b",x"fb",x"d9",x"c2"),
   576 => (x"8a",x"c2",x"4a",x"73"),
   577 => (x"bf",x"ce",x"d5",x"c2"),
   578 => (x"d9",x"c2",x"92",x"49"),
   579 => (x"72",x"48",x"bf",x"e7"),
   580 => (x"ff",x"d9",x"c2",x"80"),
   581 => (x"c4",x"48",x"71",x"58"),
   582 => (x"de",x"d5",x"c2",x"30"),
   583 => (x"87",x"ed",x"c0",x"58"),
   584 => (x"48",x"f7",x"d9",x"c2"),
   585 => (x"bf",x"eb",x"d9",x"c2"),
   586 => (x"fb",x"d9",x"c2",x"78"),
   587 => (x"ef",x"d9",x"c2",x"48"),
   588 => (x"d5",x"c2",x"78",x"bf"),
   589 => (x"c9",x"02",x"bf",x"d6"),
   590 => (x"ce",x"d5",x"c2",x"87"),
   591 => (x"31",x"c4",x"49",x"bf"),
   592 => (x"d9",x"c2",x"87",x"c7"),
   593 => (x"c4",x"49",x"bf",x"f3"),
   594 => (x"de",x"d5",x"c2",x"31"),
   595 => (x"87",x"ec",x"f6",x"59"),
   596 => (x"5c",x"5b",x"5e",x"0e"),
   597 => (x"c0",x"4a",x"71",x"0e"),
   598 => (x"02",x"9a",x"72",x"4b"),
   599 => (x"da",x"87",x"e0",x"c0"),
   600 => (x"69",x"9f",x"49",x"a2"),
   601 => (x"d6",x"d5",x"c2",x"4b"),
   602 => (x"87",x"cf",x"02",x"bf"),
   603 => (x"9f",x"49",x"a2",x"d4"),
   604 => (x"c0",x"4c",x"49",x"69"),
   605 => (x"d0",x"9c",x"ff",x"ff"),
   606 => (x"c0",x"87",x"c2",x"34"),
   607 => (x"73",x"b3",x"74",x"4c"),
   608 => (x"87",x"ee",x"fd",x"49"),
   609 => (x"0e",x"87",x"f3",x"f5"),
   610 => (x"5d",x"5c",x"5b",x"5e"),
   611 => (x"71",x"86",x"f4",x"0e"),
   612 => (x"72",x"7e",x"c0",x"4a"),
   613 => (x"87",x"d8",x"02",x"9a"),
   614 => (x"48",x"ca",x"cd",x"c2"),
   615 => (x"cd",x"c2",x"78",x"c0"),
   616 => (x"d9",x"c2",x"48",x"c2"),
   617 => (x"c2",x"78",x"bf",x"fb"),
   618 => (x"c2",x"48",x"c6",x"cd"),
   619 => (x"78",x"bf",x"f7",x"d9"),
   620 => (x"48",x"eb",x"d5",x"c2"),
   621 => (x"d5",x"c2",x"50",x"c0"),
   622 => (x"c2",x"49",x"bf",x"da"),
   623 => (x"4a",x"bf",x"ca",x"cd"),
   624 => (x"c4",x"03",x"aa",x"71"),
   625 => (x"49",x"72",x"87",x"c9"),
   626 => (x"c0",x"05",x"99",x"cf"),
   627 => (x"ed",x"c0",x"87",x"e9"),
   628 => (x"cd",x"c2",x"48",x"de"),
   629 => (x"c2",x"78",x"bf",x"c2"),
   630 => (x"c2",x"1e",x"ce",x"cd"),
   631 => (x"49",x"bf",x"c2",x"cd"),
   632 => (x"48",x"c2",x"cd",x"c2"),
   633 => (x"71",x"78",x"a1",x"c1"),
   634 => (x"c4",x"87",x"dd",x"e6"),
   635 => (x"da",x"ed",x"c0",x"86"),
   636 => (x"ce",x"cd",x"c2",x"48"),
   637 => (x"c0",x"87",x"cc",x"78"),
   638 => (x"48",x"bf",x"da",x"ed"),
   639 => (x"c0",x"80",x"e0",x"c0"),
   640 => (x"c2",x"58",x"de",x"ed"),
   641 => (x"48",x"bf",x"ca",x"cd"),
   642 => (x"cd",x"c2",x"80",x"c1"),
   643 => (x"5a",x"27",x"58",x"ce"),
   644 => (x"bf",x"00",x"00",x"0b"),
   645 => (x"9d",x"4d",x"bf",x"97"),
   646 => (x"87",x"e3",x"c2",x"02"),
   647 => (x"02",x"ad",x"e5",x"c3"),
   648 => (x"c0",x"87",x"dc",x"c2"),
   649 => (x"4b",x"bf",x"da",x"ed"),
   650 => (x"11",x"49",x"a3",x"cb"),
   651 => (x"05",x"ac",x"cf",x"4c"),
   652 => (x"75",x"87",x"d2",x"c1"),
   653 => (x"c1",x"99",x"df",x"49"),
   654 => (x"c2",x"91",x"cd",x"89"),
   655 => (x"c1",x"81",x"de",x"d5"),
   656 => (x"51",x"12",x"4a",x"a3"),
   657 => (x"12",x"4a",x"a3",x"c3"),
   658 => (x"4a",x"a3",x"c5",x"51"),
   659 => (x"a3",x"c7",x"51",x"12"),
   660 => (x"c9",x"51",x"12",x"4a"),
   661 => (x"51",x"12",x"4a",x"a3"),
   662 => (x"12",x"4a",x"a3",x"ce"),
   663 => (x"4a",x"a3",x"d0",x"51"),
   664 => (x"a3",x"d2",x"51",x"12"),
   665 => (x"d4",x"51",x"12",x"4a"),
   666 => (x"51",x"12",x"4a",x"a3"),
   667 => (x"12",x"4a",x"a3",x"d6"),
   668 => (x"4a",x"a3",x"d8",x"51"),
   669 => (x"a3",x"dc",x"51",x"12"),
   670 => (x"de",x"51",x"12",x"4a"),
   671 => (x"51",x"12",x"4a",x"a3"),
   672 => (x"fa",x"c0",x"7e",x"c1"),
   673 => (x"c8",x"49",x"74",x"87"),
   674 => (x"eb",x"c0",x"05",x"99"),
   675 => (x"d0",x"49",x"74",x"87"),
   676 => (x"87",x"d1",x"05",x"99"),
   677 => (x"c0",x"02",x"66",x"dc"),
   678 => (x"49",x"73",x"87",x"cb"),
   679 => (x"70",x"0f",x"66",x"dc"),
   680 => (x"d3",x"c0",x"02",x"98"),
   681 => (x"c0",x"05",x"6e",x"87"),
   682 => (x"d5",x"c2",x"87",x"c6"),
   683 => (x"50",x"c0",x"48",x"de"),
   684 => (x"bf",x"da",x"ed",x"c0"),
   685 => (x"87",x"dd",x"c2",x"48"),
   686 => (x"48",x"eb",x"d5",x"c2"),
   687 => (x"c2",x"7e",x"50",x"c0"),
   688 => (x"49",x"bf",x"da",x"d5"),
   689 => (x"bf",x"ca",x"cd",x"c2"),
   690 => (x"04",x"aa",x"71",x"4a"),
   691 => (x"c2",x"87",x"f7",x"fb"),
   692 => (x"05",x"bf",x"fb",x"d9"),
   693 => (x"c2",x"87",x"c8",x"c0"),
   694 => (x"02",x"bf",x"d6",x"d5"),
   695 => (x"c2",x"87",x"f4",x"c1"),
   696 => (x"49",x"bf",x"c6",x"cd"),
   697 => (x"c2",x"87",x"d9",x"f0"),
   698 => (x"c4",x"58",x"ca",x"cd"),
   699 => (x"cd",x"c2",x"48",x"a6"),
   700 => (x"c2",x"78",x"bf",x"c6"),
   701 => (x"02",x"bf",x"d6",x"d5"),
   702 => (x"c4",x"87",x"d8",x"c0"),
   703 => (x"ff",x"cf",x"49",x"66"),
   704 => (x"99",x"f8",x"ff",x"ff"),
   705 => (x"c5",x"c0",x"02",x"a9"),
   706 => (x"c0",x"4c",x"c0",x"87"),
   707 => (x"4c",x"c1",x"87",x"e1"),
   708 => (x"c4",x"87",x"dc",x"c0"),
   709 => (x"ff",x"cf",x"49",x"66"),
   710 => (x"02",x"a9",x"99",x"f8"),
   711 => (x"c8",x"87",x"c8",x"c0"),
   712 => (x"78",x"c0",x"48",x"a6"),
   713 => (x"c8",x"87",x"c5",x"c0"),
   714 => (x"78",x"c1",x"48",x"a6"),
   715 => (x"74",x"4c",x"66",x"c8"),
   716 => (x"de",x"c0",x"05",x"9c"),
   717 => (x"49",x"66",x"c4",x"87"),
   718 => (x"d5",x"c2",x"89",x"c2"),
   719 => (x"c2",x"91",x"bf",x"ce"),
   720 => (x"48",x"bf",x"e7",x"d9"),
   721 => (x"cd",x"c2",x"80",x"71"),
   722 => (x"cd",x"c2",x"58",x"c6"),
   723 => (x"78",x"c0",x"48",x"ca"),
   724 => (x"c0",x"87",x"e3",x"f9"),
   725 => (x"ee",x"8e",x"f4",x"48"),
   726 => (x"00",x"00",x"87",x"de"),
   727 => (x"ff",x"ff",x"00",x"00"),
   728 => (x"0b",x"6a",x"ff",x"ff"),
   729 => (x"0b",x"73",x"00",x"00"),
   730 => (x"41",x"46",x"00",x"00"),
   731 => (x"20",x"32",x"33",x"54"),
   732 => (x"46",x"00",x"20",x"20"),
   733 => (x"36",x"31",x"54",x"41"),
   734 => (x"00",x"20",x"20",x"20"),
   735 => (x"48",x"d4",x"ff",x"1e"),
   736 => (x"68",x"78",x"ff",x"c3"),
   737 => (x"1e",x"4f",x"26",x"48"),
   738 => (x"c3",x"48",x"d4",x"ff"),
   739 => (x"d0",x"ff",x"78",x"ff"),
   740 => (x"78",x"e1",x"c0",x"48"),
   741 => (x"d4",x"48",x"d4",x"ff"),
   742 => (x"ff",x"d9",x"c2",x"78"),
   743 => (x"bf",x"d4",x"ff",x"48"),
   744 => (x"1e",x"4f",x"26",x"50"),
   745 => (x"c0",x"48",x"d0",x"ff"),
   746 => (x"4f",x"26",x"78",x"e0"),
   747 => (x"87",x"cc",x"ff",x"1e"),
   748 => (x"02",x"99",x"49",x"70"),
   749 => (x"fb",x"c0",x"87",x"c6"),
   750 => (x"87",x"f1",x"05",x"a9"),
   751 => (x"4f",x"26",x"48",x"71"),
   752 => (x"5c",x"5b",x"5e",x"0e"),
   753 => (x"c0",x"4b",x"71",x"0e"),
   754 => (x"87",x"f0",x"fe",x"4c"),
   755 => (x"02",x"99",x"49",x"70"),
   756 => (x"c0",x"87",x"f9",x"c0"),
   757 => (x"c0",x"02",x"a9",x"ec"),
   758 => (x"fb",x"c0",x"87",x"f2"),
   759 => (x"eb",x"c0",x"02",x"a9"),
   760 => (x"b7",x"66",x"cc",x"87"),
   761 => (x"87",x"c7",x"03",x"ac"),
   762 => (x"c2",x"02",x"66",x"d0"),
   763 => (x"71",x"53",x"71",x"87"),
   764 => (x"87",x"c2",x"02",x"99"),
   765 => (x"c3",x"fe",x"84",x"c1"),
   766 => (x"99",x"49",x"70",x"87"),
   767 => (x"c0",x"87",x"cd",x"02"),
   768 => (x"c7",x"02",x"a9",x"ec"),
   769 => (x"a9",x"fb",x"c0",x"87"),
   770 => (x"87",x"d5",x"ff",x"05"),
   771 => (x"c3",x"02",x"66",x"d0"),
   772 => (x"7b",x"97",x"c0",x"87"),
   773 => (x"05",x"a9",x"ec",x"c0"),
   774 => (x"4a",x"74",x"87",x"c4"),
   775 => (x"4a",x"74",x"87",x"c5"),
   776 => (x"72",x"8a",x"0a",x"c0"),
   777 => (x"26",x"87",x"c2",x"48"),
   778 => (x"26",x"4c",x"26",x"4d"),
   779 => (x"1e",x"4f",x"26",x"4b"),
   780 => (x"70",x"87",x"c9",x"fd"),
   781 => (x"a9",x"f0",x"c0",x"49"),
   782 => (x"c0",x"87",x"c9",x"04"),
   783 => (x"c3",x"01",x"a9",x"f9"),
   784 => (x"89",x"f0",x"c0",x"87"),
   785 => (x"04",x"a9",x"c1",x"c1"),
   786 => (x"da",x"c1",x"87",x"c9"),
   787 => (x"87",x"c3",x"01",x"a9"),
   788 => (x"71",x"89",x"f7",x"c0"),
   789 => (x"0e",x"4f",x"26",x"48"),
   790 => (x"5d",x"5c",x"5b",x"5e"),
   791 => (x"71",x"86",x"f8",x"0e"),
   792 => (x"fc",x"4d",x"c0",x"4c"),
   793 => (x"4b",x"c0",x"87",x"e1"),
   794 => (x"97",x"f6",x"f3",x"c0"),
   795 => (x"a9",x"c0",x"49",x"bf"),
   796 => (x"fc",x"87",x"cf",x"04"),
   797 => (x"83",x"c1",x"87",x"f6"),
   798 => (x"97",x"f6",x"f3",x"c0"),
   799 => (x"06",x"ab",x"49",x"bf"),
   800 => (x"f3",x"c0",x"87",x"f1"),
   801 => (x"02",x"bf",x"97",x"f6"),
   802 => (x"ef",x"fb",x"87",x"cf"),
   803 => (x"99",x"49",x"70",x"87"),
   804 => (x"c0",x"87",x"c6",x"02"),
   805 => (x"f1",x"05",x"a9",x"ec"),
   806 => (x"fb",x"4b",x"c0",x"87"),
   807 => (x"7e",x"70",x"87",x"de"),
   808 => (x"c8",x"87",x"d9",x"fb"),
   809 => (x"d3",x"fb",x"58",x"a6"),
   810 => (x"c1",x"4a",x"70",x"87"),
   811 => (x"49",x"a4",x"c8",x"83"),
   812 => (x"6e",x"49",x"69",x"97"),
   813 => (x"87",x"da",x"05",x"a9"),
   814 => (x"97",x"49",x"a4",x"c9"),
   815 => (x"66",x"c4",x"49",x"69"),
   816 => (x"87",x"ce",x"05",x"a9"),
   817 => (x"97",x"49",x"a4",x"ca"),
   818 => (x"05",x"aa",x"49",x"69"),
   819 => (x"4d",x"c1",x"87",x"c4"),
   820 => (x"48",x"6e",x"87",x"d4"),
   821 => (x"02",x"a8",x"ec",x"c0"),
   822 => (x"48",x"6e",x"87",x"c8"),
   823 => (x"05",x"a8",x"fb",x"c0"),
   824 => (x"4b",x"c0",x"87",x"c4"),
   825 => (x"9d",x"75",x"4d",x"c1"),
   826 => (x"87",x"ef",x"fe",x"02"),
   827 => (x"73",x"87",x"f4",x"fa"),
   828 => (x"fc",x"8e",x"f8",x"48"),
   829 => (x"0e",x"00",x"87",x"f1"),
   830 => (x"5d",x"5c",x"5b",x"5e"),
   831 => (x"71",x"86",x"f8",x"0e"),
   832 => (x"4b",x"d4",x"ff",x"7e"),
   833 => (x"da",x"c2",x"1e",x"6e"),
   834 => (x"e5",x"e9",x"49",x"c4"),
   835 => (x"70",x"86",x"c4",x"87"),
   836 => (x"ea",x"c4",x"02",x"98"),
   837 => (x"dd",x"dd",x"c1",x"87"),
   838 => (x"49",x"6e",x"4d",x"bf"),
   839 => (x"c8",x"87",x"f8",x"fc"),
   840 => (x"98",x"70",x"58",x"a6"),
   841 => (x"c4",x"87",x"c5",x"05"),
   842 => (x"78",x"c1",x"48",x"a6"),
   843 => (x"c5",x"48",x"d0",x"ff"),
   844 => (x"7b",x"d5",x"c1",x"78"),
   845 => (x"c1",x"49",x"66",x"c4"),
   846 => (x"c1",x"31",x"c6",x"89"),
   847 => (x"bf",x"97",x"db",x"dd"),
   848 => (x"b0",x"71",x"48",x"4a"),
   849 => (x"d0",x"ff",x"7b",x"70"),
   850 => (x"c2",x"78",x"c4",x"48"),
   851 => (x"bf",x"97",x"ff",x"d9"),
   852 => (x"02",x"99",x"d0",x"49"),
   853 => (x"78",x"c5",x"87",x"d7"),
   854 => (x"c0",x"7b",x"d6",x"c1"),
   855 => (x"7b",x"ff",x"c3",x"4a"),
   856 => (x"e0",x"c0",x"82",x"c1"),
   857 => (x"87",x"f5",x"04",x"aa"),
   858 => (x"c4",x"48",x"d0",x"ff"),
   859 => (x"7b",x"ff",x"c3",x"78"),
   860 => (x"c5",x"48",x"d0",x"ff"),
   861 => (x"7b",x"d3",x"c1",x"78"),
   862 => (x"78",x"c4",x"7b",x"c1"),
   863 => (x"06",x"ad",x"b7",x"c0"),
   864 => (x"c2",x"87",x"eb",x"c2"),
   865 => (x"4c",x"bf",x"cc",x"da"),
   866 => (x"c2",x"02",x"9c",x"8d"),
   867 => (x"cd",x"c2",x"87",x"c2"),
   868 => (x"a6",x"c4",x"7e",x"ce"),
   869 => (x"78",x"c0",x"c8",x"48"),
   870 => (x"ac",x"b7",x"c0",x"8c"),
   871 => (x"c8",x"87",x"c6",x"03"),
   872 => (x"c0",x"78",x"a4",x"c0"),
   873 => (x"ff",x"d9",x"c2",x"4c"),
   874 => (x"d0",x"49",x"bf",x"97"),
   875 => (x"87",x"d0",x"02",x"99"),
   876 => (x"da",x"c2",x"1e",x"c0"),
   877 => (x"eb",x"eb",x"49",x"c4"),
   878 => (x"70",x"86",x"c4",x"87"),
   879 => (x"87",x"f5",x"c0",x"4a"),
   880 => (x"1e",x"ce",x"cd",x"c2"),
   881 => (x"49",x"c4",x"da",x"c2"),
   882 => (x"c4",x"87",x"d9",x"eb"),
   883 => (x"ff",x"4a",x"70",x"86"),
   884 => (x"c5",x"c8",x"48",x"d0"),
   885 => (x"7b",x"d4",x"c1",x"78"),
   886 => (x"7b",x"bf",x"97",x"6e"),
   887 => (x"80",x"c1",x"48",x"6e"),
   888 => (x"66",x"c4",x"7e",x"70"),
   889 => (x"c8",x"88",x"c1",x"48"),
   890 => (x"98",x"70",x"58",x"a6"),
   891 => (x"87",x"e8",x"ff",x"05"),
   892 => (x"c4",x"48",x"d0",x"ff"),
   893 => (x"05",x"9a",x"72",x"78"),
   894 => (x"48",x"c0",x"87",x"c5"),
   895 => (x"c1",x"87",x"c2",x"c1"),
   896 => (x"c4",x"da",x"c2",x"1e"),
   897 => (x"87",x"c2",x"e9",x"49"),
   898 => (x"9c",x"74",x"86",x"c4"),
   899 => (x"87",x"fe",x"fd",x"05"),
   900 => (x"06",x"ad",x"b7",x"c0"),
   901 => (x"da",x"c2",x"87",x"d1"),
   902 => (x"78",x"c0",x"48",x"c4"),
   903 => (x"78",x"c0",x"80",x"d0"),
   904 => (x"da",x"c2",x"80",x"f4"),
   905 => (x"c0",x"78",x"bf",x"d0"),
   906 => (x"fd",x"01",x"ad",x"b7"),
   907 => (x"d0",x"ff",x"87",x"d5"),
   908 => (x"c1",x"78",x"c5",x"48"),
   909 => (x"7b",x"c0",x"7b",x"d3"),
   910 => (x"48",x"c1",x"78",x"c4"),
   911 => (x"c0",x"87",x"c2",x"c0"),
   912 => (x"26",x"8e",x"f8",x"48"),
   913 => (x"26",x"4c",x"26",x"4d"),
   914 => (x"0e",x"4f",x"26",x"4b"),
   915 => (x"5d",x"5c",x"5b",x"5e"),
   916 => (x"4b",x"71",x"1e",x"0e"),
   917 => (x"ab",x"4d",x"4c",x"c0"),
   918 => (x"87",x"e8",x"c0",x"04"),
   919 => (x"1e",x"d7",x"f1",x"c0"),
   920 => (x"c4",x"02",x"9d",x"75"),
   921 => (x"c2",x"4a",x"c0",x"87"),
   922 => (x"72",x"4a",x"c1",x"87"),
   923 => (x"87",x"d7",x"ec",x"49"),
   924 => (x"7e",x"70",x"86",x"c4"),
   925 => (x"05",x"6e",x"84",x"c1"),
   926 => (x"4c",x"73",x"87",x"c2"),
   927 => (x"ac",x"73",x"85",x"c1"),
   928 => (x"87",x"d8",x"ff",x"06"),
   929 => (x"fe",x"26",x"48",x"6e"),
   930 => (x"71",x"1e",x"87",x"f9"),
   931 => (x"05",x"66",x"c4",x"4a"),
   932 => (x"49",x"72",x"87",x"c5"),
   933 => (x"26",x"87",x"e0",x"f9"),
   934 => (x"5b",x"5e",x"0e",x"4f"),
   935 => (x"1e",x"0e",x"5d",x"5c"),
   936 => (x"de",x"49",x"4c",x"71"),
   937 => (x"ec",x"da",x"c2",x"91"),
   938 => (x"97",x"85",x"71",x"4d"),
   939 => (x"dc",x"c1",x"02",x"6d"),
   940 => (x"d8",x"da",x"c2",x"87"),
   941 => (x"81",x"74",x"49",x"bf"),
   942 => (x"87",x"cf",x"fe",x"71"),
   943 => (x"98",x"48",x"7e",x"70"),
   944 => (x"87",x"f2",x"c0",x"02"),
   945 => (x"4b",x"e0",x"da",x"c2"),
   946 => (x"49",x"cb",x"4a",x"70"),
   947 => (x"87",x"d7",x"c7",x"ff"),
   948 => (x"93",x"cb",x"4b",x"74"),
   949 => (x"83",x"ef",x"dd",x"c1"),
   950 => (x"fc",x"c0",x"83",x"c4"),
   951 => (x"49",x"74",x"7b",x"d1"),
   952 => (x"87",x"e9",x"c0",x"c1"),
   953 => (x"dd",x"c1",x"7b",x"75"),
   954 => (x"49",x"bf",x"97",x"dc"),
   955 => (x"e0",x"da",x"c2",x"1e"),
   956 => (x"87",x"d6",x"fe",x"49"),
   957 => (x"49",x"74",x"86",x"c4"),
   958 => (x"87",x"d1",x"c0",x"c1"),
   959 => (x"c1",x"c1",x"49",x"c0"),
   960 => (x"da",x"c2",x"87",x"f0"),
   961 => (x"78",x"c0",x"48",x"c0"),
   962 => (x"f9",x"dd",x"49",x"c1"),
   963 => (x"f2",x"fc",x"26",x"87"),
   964 => (x"61",x"6f",x"4c",x"87"),
   965 => (x"67",x"6e",x"69",x"64"),
   966 => (x"00",x"2e",x"2e",x"2e"),
   967 => (x"71",x"1e",x"73",x"1e"),
   968 => (x"da",x"c2",x"49",x"4a"),
   969 => (x"71",x"81",x"bf",x"d8"),
   970 => (x"70",x"87",x"e0",x"fc"),
   971 => (x"c4",x"02",x"9b",x"4b"),
   972 => (x"db",x"e8",x"49",x"87"),
   973 => (x"d8",x"da",x"c2",x"87"),
   974 => (x"c1",x"78",x"c0",x"48"),
   975 => (x"87",x"c6",x"dd",x"49"),
   976 => (x"1e",x"87",x"c4",x"fc"),
   977 => (x"c0",x"c1",x"49",x"c0"),
   978 => (x"4f",x"26",x"87",x"e8"),
   979 => (x"49",x"4a",x"71",x"1e"),
   980 => (x"dd",x"c1",x"91",x"cb"),
   981 => (x"81",x"c8",x"81",x"ef"),
   982 => (x"da",x"c2",x"48",x"11"),
   983 => (x"da",x"c2",x"58",x"c4"),
   984 => (x"78",x"c0",x"48",x"d8"),
   985 => (x"dd",x"dc",x"49",x"c1"),
   986 => (x"1e",x"4f",x"26",x"87"),
   987 => (x"d2",x"02",x"99",x"71"),
   988 => (x"c4",x"df",x"c1",x"87"),
   989 => (x"f7",x"50",x"c0",x"48"),
   990 => (x"cc",x"fd",x"c0",x"80"),
   991 => (x"e8",x"dd",x"c1",x"40"),
   992 => (x"c1",x"87",x"ce",x"78"),
   993 => (x"c1",x"48",x"c0",x"df"),
   994 => (x"fc",x"78",x"e1",x"dd"),
   995 => (x"c3",x"fd",x"c0",x"80"),
   996 => (x"0e",x"4f",x"26",x"78"),
   997 => (x"5d",x"5c",x"5b",x"5e"),
   998 => (x"c2",x"86",x"f4",x"0e"),
   999 => (x"c0",x"4d",x"ce",x"cd"),
  1000 => (x"48",x"a6",x"c4",x"4c"),
  1001 => (x"da",x"c2",x"78",x"c0"),
  1002 => (x"c0",x"48",x"bf",x"d8"),
  1003 => (x"c0",x"c1",x"06",x"a8"),
  1004 => (x"ce",x"cd",x"c2",x"87"),
  1005 => (x"c0",x"02",x"98",x"48"),
  1006 => (x"f1",x"c0",x"87",x"f7"),
  1007 => (x"66",x"c8",x"1e",x"d7"),
  1008 => (x"c4",x"87",x"c7",x"02"),
  1009 => (x"78",x"c0",x"48",x"a6"),
  1010 => (x"a6",x"c4",x"87",x"c5"),
  1011 => (x"c4",x"78",x"c1",x"48"),
  1012 => (x"f2",x"e6",x"49",x"66"),
  1013 => (x"70",x"86",x"c4",x"87"),
  1014 => (x"c4",x"84",x"c1",x"4d"),
  1015 => (x"80",x"c1",x"48",x"66"),
  1016 => (x"c2",x"58",x"a6",x"c8"),
  1017 => (x"ac",x"bf",x"d8",x"da"),
  1018 => (x"75",x"87",x"c6",x"03"),
  1019 => (x"c9",x"ff",x"05",x"9d"),
  1020 => (x"75",x"4c",x"c0",x"87"),
  1021 => (x"dc",x"c3",x"02",x"9d"),
  1022 => (x"d7",x"f1",x"c0",x"87"),
  1023 => (x"02",x"66",x"c8",x"1e"),
  1024 => (x"a6",x"cc",x"87",x"c7"),
  1025 => (x"c5",x"78",x"c0",x"48"),
  1026 => (x"48",x"a6",x"cc",x"87"),
  1027 => (x"66",x"cc",x"78",x"c1"),
  1028 => (x"87",x"f3",x"e5",x"49"),
  1029 => (x"7e",x"70",x"86",x"c4"),
  1030 => (x"c2",x"02",x"98",x"48"),
  1031 => (x"cb",x"49",x"87",x"e4"),
  1032 => (x"49",x"69",x"97",x"81"),
  1033 => (x"c1",x"02",x"99",x"d0"),
  1034 => (x"49",x"74",x"87",x"d4"),
  1035 => (x"dd",x"c1",x"91",x"cb"),
  1036 => (x"fc",x"c0",x"81",x"ef"),
  1037 => (x"81",x"c8",x"79",x"dc"),
  1038 => (x"74",x"51",x"ff",x"c3"),
  1039 => (x"c2",x"91",x"de",x"49"),
  1040 => (x"71",x"4d",x"ec",x"da"),
  1041 => (x"97",x"c1",x"c2",x"85"),
  1042 => (x"49",x"a5",x"c1",x"7d"),
  1043 => (x"c2",x"51",x"e0",x"c0"),
  1044 => (x"bf",x"97",x"de",x"d5"),
  1045 => (x"c1",x"87",x"d2",x"02"),
  1046 => (x"4b",x"a5",x"c2",x"84"),
  1047 => (x"4a",x"de",x"d5",x"c2"),
  1048 => (x"c1",x"ff",x"49",x"db"),
  1049 => (x"d9",x"c1",x"87",x"c1"),
  1050 => (x"49",x"a5",x"cd",x"87"),
  1051 => (x"84",x"c1",x"51",x"c0"),
  1052 => (x"6e",x"4b",x"a5",x"c2"),
  1053 => (x"ff",x"49",x"cb",x"4a"),
  1054 => (x"c1",x"87",x"ec",x"c0"),
  1055 => (x"49",x"74",x"87",x"c4"),
  1056 => (x"dd",x"c1",x"91",x"cb"),
  1057 => (x"fa",x"c0",x"81",x"ef"),
  1058 => (x"d5",x"c2",x"79",x"d9"),
  1059 => (x"02",x"bf",x"97",x"de"),
  1060 => (x"49",x"74",x"87",x"d8"),
  1061 => (x"84",x"c1",x"91",x"de"),
  1062 => (x"4b",x"ec",x"da",x"c2"),
  1063 => (x"d5",x"c2",x"83",x"71"),
  1064 => (x"49",x"dd",x"4a",x"de"),
  1065 => (x"87",x"ff",x"ff",x"fe"),
  1066 => (x"4b",x"74",x"87",x"d8"),
  1067 => (x"da",x"c2",x"93",x"de"),
  1068 => (x"a3",x"cb",x"83",x"ec"),
  1069 => (x"c1",x"51",x"c0",x"49"),
  1070 => (x"4a",x"6e",x"73",x"84"),
  1071 => (x"ff",x"fe",x"49",x"cb"),
  1072 => (x"66",x"c4",x"87",x"e5"),
  1073 => (x"c8",x"80",x"c1",x"48"),
  1074 => (x"ac",x"c7",x"58",x"a6"),
  1075 => (x"87",x"c5",x"c0",x"03"),
  1076 => (x"e4",x"fc",x"05",x"6e"),
  1077 => (x"f4",x"48",x"74",x"87"),
  1078 => (x"87",x"e7",x"f5",x"8e"),
  1079 => (x"71",x"1e",x"73",x"1e"),
  1080 => (x"91",x"cb",x"49",x"4b"),
  1081 => (x"81",x"ef",x"dd",x"c1"),
  1082 => (x"c1",x"4a",x"a1",x"c8"),
  1083 => (x"12",x"48",x"db",x"dd"),
  1084 => (x"4a",x"a1",x"c9",x"50"),
  1085 => (x"48",x"f6",x"f3",x"c0"),
  1086 => (x"81",x"ca",x"50",x"12"),
  1087 => (x"48",x"dc",x"dd",x"c1"),
  1088 => (x"dd",x"c1",x"50",x"11"),
  1089 => (x"49",x"bf",x"97",x"dc"),
  1090 => (x"f5",x"49",x"c0",x"1e"),
  1091 => (x"da",x"c2",x"87",x"fc"),
  1092 => (x"78",x"de",x"48",x"c0"),
  1093 => (x"ed",x"d5",x"49",x"c1"),
  1094 => (x"ea",x"f4",x"26",x"87"),
  1095 => (x"5b",x"5e",x"0e",x"87"),
  1096 => (x"f4",x"0e",x"5d",x"5c"),
  1097 => (x"49",x"4d",x"71",x"86"),
  1098 => (x"dd",x"c1",x"91",x"cb"),
  1099 => (x"a1",x"c8",x"81",x"ef"),
  1100 => (x"7e",x"a1",x"ca",x"4a"),
  1101 => (x"c2",x"48",x"a6",x"c4"),
  1102 => (x"78",x"bf",x"c8",x"de"),
  1103 => (x"4b",x"bf",x"97",x"6e"),
  1104 => (x"73",x"4c",x"66",x"c4"),
  1105 => (x"cc",x"48",x"12",x"2c"),
  1106 => (x"9c",x"70",x"58",x"a6"),
  1107 => (x"81",x"c9",x"84",x"c1"),
  1108 => (x"b7",x"49",x"69",x"97"),
  1109 => (x"87",x"c2",x"04",x"ac"),
  1110 => (x"97",x"6e",x"4c",x"c0"),
  1111 => (x"66",x"c8",x"4a",x"bf"),
  1112 => (x"ff",x"31",x"72",x"49"),
  1113 => (x"99",x"66",x"c4",x"b9"),
  1114 => (x"30",x"72",x"48",x"74"),
  1115 => (x"71",x"48",x"4a",x"70"),
  1116 => (x"cc",x"de",x"c2",x"b0"),
  1117 => (x"d4",x"e4",x"c0",x"58"),
  1118 => (x"d4",x"49",x"c0",x"87"),
  1119 => (x"49",x"75",x"87",x"c8"),
  1120 => (x"87",x"c9",x"f6",x"c0"),
  1121 => (x"fa",x"f2",x"8e",x"f4"),
  1122 => (x"1e",x"73",x"1e",x"87"),
  1123 => (x"fe",x"49",x"4b",x"71"),
  1124 => (x"49",x"73",x"87",x"cb"),
  1125 => (x"f2",x"87",x"c6",x"fe"),
  1126 => (x"73",x"1e",x"87",x"ed"),
  1127 => (x"c6",x"4b",x"71",x"1e"),
  1128 => (x"db",x"02",x"4a",x"a3"),
  1129 => (x"02",x"8a",x"c1",x"87"),
  1130 => (x"02",x"8a",x"87",x"d6"),
  1131 => (x"8a",x"87",x"da",x"c1"),
  1132 => (x"87",x"fc",x"c0",x"02"),
  1133 => (x"e1",x"c0",x"02",x"8a"),
  1134 => (x"cb",x"02",x"8a",x"87"),
  1135 => (x"87",x"db",x"c1",x"87"),
  1136 => (x"c7",x"f6",x"49",x"c7"),
  1137 => (x"87",x"de",x"c1",x"87"),
  1138 => (x"bf",x"d8",x"da",x"c2"),
  1139 => (x"87",x"cb",x"c1",x"02"),
  1140 => (x"c2",x"88",x"c1",x"48"),
  1141 => (x"c1",x"58",x"dc",x"da"),
  1142 => (x"da",x"c2",x"87",x"c1"),
  1143 => (x"c0",x"02",x"bf",x"dc"),
  1144 => (x"da",x"c2",x"87",x"f9"),
  1145 => (x"c1",x"48",x"bf",x"d8"),
  1146 => (x"dc",x"da",x"c2",x"80"),
  1147 => (x"87",x"eb",x"c0",x"58"),
  1148 => (x"bf",x"d8",x"da",x"c2"),
  1149 => (x"c2",x"89",x"c6",x"49"),
  1150 => (x"c0",x"59",x"dc",x"da"),
  1151 => (x"da",x"03",x"a9",x"b7"),
  1152 => (x"d8",x"da",x"c2",x"87"),
  1153 => (x"d2",x"78",x"c0",x"48"),
  1154 => (x"dc",x"da",x"c2",x"87"),
  1155 => (x"87",x"cb",x"02",x"bf"),
  1156 => (x"bf",x"d8",x"da",x"c2"),
  1157 => (x"c2",x"80",x"c6",x"48"),
  1158 => (x"c0",x"58",x"dc",x"da"),
  1159 => (x"87",x"e6",x"d1",x"49"),
  1160 => (x"f3",x"c0",x"49",x"73"),
  1161 => (x"de",x"f0",x"87",x"e7"),
  1162 => (x"5b",x"5e",x"0e",x"87"),
  1163 => (x"ff",x"0e",x"5d",x"5c"),
  1164 => (x"a6",x"dc",x"86",x"d4"),
  1165 => (x"48",x"a6",x"c8",x"59"),
  1166 => (x"80",x"c4",x"78",x"c0"),
  1167 => (x"78",x"66",x"c0",x"c1"),
  1168 => (x"78",x"c1",x"80",x"c4"),
  1169 => (x"78",x"c1",x"80",x"c4"),
  1170 => (x"48",x"dc",x"da",x"c2"),
  1171 => (x"da",x"c2",x"78",x"c1"),
  1172 => (x"de",x"48",x"bf",x"c0"),
  1173 => (x"87",x"c9",x"05",x"a8"),
  1174 => (x"cc",x"87",x"f8",x"f4"),
  1175 => (x"e4",x"cf",x"58",x"a6"),
  1176 => (x"87",x"e3",x"e4",x"87"),
  1177 => (x"e4",x"87",x"c5",x"e5"),
  1178 => (x"4c",x"70",x"87",x"d2"),
  1179 => (x"02",x"ac",x"fb",x"c0"),
  1180 => (x"d8",x"87",x"fb",x"c1"),
  1181 => (x"ed",x"c1",x"05",x"66"),
  1182 => (x"66",x"fc",x"c0",x"87"),
  1183 => (x"6a",x"82",x"c4",x"4a"),
  1184 => (x"c1",x"1e",x"72",x"7e"),
  1185 => (x"c4",x"48",x"fa",x"d9"),
  1186 => (x"a1",x"c8",x"49",x"66"),
  1187 => (x"71",x"41",x"20",x"4a"),
  1188 => (x"87",x"f9",x"05",x"aa"),
  1189 => (x"4a",x"26",x"51",x"10"),
  1190 => (x"48",x"66",x"fc",x"c0"),
  1191 => (x"78",x"dc",x"c3",x"c1"),
  1192 => (x"81",x"c7",x"49",x"6a"),
  1193 => (x"fc",x"c0",x"51",x"74"),
  1194 => (x"81",x"c8",x"49",x"66"),
  1195 => (x"fc",x"c0",x"51",x"c1"),
  1196 => (x"81",x"c9",x"49",x"66"),
  1197 => (x"fc",x"c0",x"51",x"c0"),
  1198 => (x"81",x"ca",x"49",x"66"),
  1199 => (x"1e",x"c1",x"51",x"c0"),
  1200 => (x"49",x"6a",x"1e",x"d8"),
  1201 => (x"f7",x"e3",x"81",x"c8"),
  1202 => (x"c1",x"86",x"c8",x"87"),
  1203 => (x"c0",x"48",x"66",x"c0"),
  1204 => (x"87",x"c7",x"01",x"a8"),
  1205 => (x"c1",x"48",x"a6",x"c8"),
  1206 => (x"c1",x"87",x"ce",x"78"),
  1207 => (x"c1",x"48",x"66",x"c0"),
  1208 => (x"58",x"a6",x"d0",x"88"),
  1209 => (x"c3",x"e3",x"87",x"c3"),
  1210 => (x"48",x"a6",x"d0",x"87"),
  1211 => (x"9c",x"74",x"78",x"c2"),
  1212 => (x"87",x"cd",x"cd",x"02"),
  1213 => (x"c1",x"48",x"66",x"c8"),
  1214 => (x"03",x"a8",x"66",x"c4"),
  1215 => (x"dc",x"87",x"c2",x"cd"),
  1216 => (x"78",x"c0",x"48",x"a6"),
  1217 => (x"78",x"c0",x"80",x"e8"),
  1218 => (x"70",x"87",x"f1",x"e1"),
  1219 => (x"ac",x"d0",x"c1",x"4c"),
  1220 => (x"87",x"d5",x"c2",x"05"),
  1221 => (x"e4",x"7e",x"66",x"c4"),
  1222 => (x"a6",x"c8",x"87",x"d5"),
  1223 => (x"87",x"dc",x"e1",x"58"),
  1224 => (x"ec",x"c0",x"4c",x"70"),
  1225 => (x"eb",x"c1",x"05",x"ac"),
  1226 => (x"49",x"66",x"c8",x"87"),
  1227 => (x"fc",x"c0",x"91",x"cb"),
  1228 => (x"a1",x"c4",x"81",x"66"),
  1229 => (x"c8",x"4d",x"6a",x"4a"),
  1230 => (x"66",x"c4",x"4a",x"a1"),
  1231 => (x"cc",x"fd",x"c0",x"52"),
  1232 => (x"87",x"f8",x"e0",x"79"),
  1233 => (x"02",x"9c",x"4c",x"70"),
  1234 => (x"fb",x"c0",x"87",x"d8"),
  1235 => (x"87",x"d2",x"02",x"ac"),
  1236 => (x"e7",x"e0",x"55",x"74"),
  1237 => (x"9c",x"4c",x"70",x"87"),
  1238 => (x"c0",x"87",x"c7",x"02"),
  1239 => (x"ff",x"05",x"ac",x"fb"),
  1240 => (x"e0",x"c0",x"87",x"ee"),
  1241 => (x"55",x"c1",x"c2",x"55"),
  1242 => (x"d8",x"7d",x"97",x"c0"),
  1243 => (x"a8",x"6e",x"48",x"66"),
  1244 => (x"c8",x"87",x"db",x"05"),
  1245 => (x"66",x"cc",x"48",x"66"),
  1246 => (x"87",x"ca",x"04",x"a8"),
  1247 => (x"c1",x"48",x"66",x"c8"),
  1248 => (x"58",x"a6",x"cc",x"80"),
  1249 => (x"66",x"cc",x"87",x"c8"),
  1250 => (x"d0",x"88",x"c1",x"48"),
  1251 => (x"df",x"ff",x"58",x"a6"),
  1252 => (x"4c",x"70",x"87",x"ea"),
  1253 => (x"05",x"ac",x"d0",x"c1"),
  1254 => (x"66",x"d4",x"87",x"c8"),
  1255 => (x"d8",x"80",x"c1",x"48"),
  1256 => (x"d0",x"c1",x"58",x"a6"),
  1257 => (x"eb",x"fd",x"02",x"ac"),
  1258 => (x"48",x"66",x"c4",x"87"),
  1259 => (x"05",x"a8",x"66",x"d8"),
  1260 => (x"c0",x"87",x"e0",x"c9"),
  1261 => (x"c0",x"48",x"a6",x"e0"),
  1262 => (x"c0",x"48",x"74",x"78"),
  1263 => (x"7e",x"70",x"88",x"fb"),
  1264 => (x"c9",x"02",x"98",x"48"),
  1265 => (x"cb",x"48",x"87",x"e2"),
  1266 => (x"48",x"7e",x"70",x"88"),
  1267 => (x"cd",x"c1",x"02",x"98"),
  1268 => (x"88",x"c9",x"48",x"87"),
  1269 => (x"98",x"48",x"7e",x"70"),
  1270 => (x"87",x"fe",x"c3",x"02"),
  1271 => (x"70",x"88",x"c4",x"48"),
  1272 => (x"02",x"98",x"48",x"7e"),
  1273 => (x"c1",x"48",x"87",x"ce"),
  1274 => (x"48",x"7e",x"70",x"88"),
  1275 => (x"e9",x"c3",x"02",x"98"),
  1276 => (x"87",x"d6",x"c8",x"87"),
  1277 => (x"c0",x"48",x"a6",x"dc"),
  1278 => (x"dd",x"ff",x"78",x"f0"),
  1279 => (x"4c",x"70",x"87",x"fe"),
  1280 => (x"02",x"ac",x"ec",x"c0"),
  1281 => (x"c0",x"87",x"c4",x"c0"),
  1282 => (x"c0",x"5c",x"a6",x"e0"),
  1283 => (x"cd",x"02",x"ac",x"ec"),
  1284 => (x"e7",x"dd",x"ff",x"87"),
  1285 => (x"c0",x"4c",x"70",x"87"),
  1286 => (x"ff",x"05",x"ac",x"ec"),
  1287 => (x"ec",x"c0",x"87",x"f3"),
  1288 => (x"c4",x"c0",x"02",x"ac"),
  1289 => (x"d3",x"dd",x"ff",x"87"),
  1290 => (x"ca",x"1e",x"c0",x"87"),
  1291 => (x"49",x"66",x"d0",x"1e"),
  1292 => (x"c4",x"c1",x"91",x"cb"),
  1293 => (x"80",x"71",x"48",x"66"),
  1294 => (x"c8",x"58",x"a6",x"cc"),
  1295 => (x"80",x"c4",x"48",x"66"),
  1296 => (x"cc",x"58",x"a6",x"d0"),
  1297 => (x"ff",x"49",x"bf",x"66"),
  1298 => (x"c1",x"87",x"f5",x"dd"),
  1299 => (x"d4",x"1e",x"de",x"1e"),
  1300 => (x"ff",x"49",x"bf",x"66"),
  1301 => (x"d0",x"87",x"e9",x"dd"),
  1302 => (x"48",x"49",x"70",x"86"),
  1303 => (x"c0",x"88",x"08",x"c0"),
  1304 => (x"c0",x"58",x"a6",x"e8"),
  1305 => (x"ee",x"c0",x"06",x"a8"),
  1306 => (x"66",x"e4",x"c0",x"87"),
  1307 => (x"03",x"a8",x"dd",x"48"),
  1308 => (x"c4",x"87",x"e4",x"c0"),
  1309 => (x"c0",x"49",x"bf",x"66"),
  1310 => (x"c0",x"81",x"66",x"e4"),
  1311 => (x"e4",x"c0",x"51",x"e0"),
  1312 => (x"81",x"c1",x"49",x"66"),
  1313 => (x"81",x"bf",x"66",x"c4"),
  1314 => (x"c0",x"51",x"c1",x"c2"),
  1315 => (x"c2",x"49",x"66",x"e4"),
  1316 => (x"bf",x"66",x"c4",x"81"),
  1317 => (x"6e",x"51",x"c0",x"81"),
  1318 => (x"dc",x"c3",x"c1",x"48"),
  1319 => (x"c8",x"49",x"6e",x"78"),
  1320 => (x"51",x"66",x"d0",x"81"),
  1321 => (x"81",x"c9",x"49",x"6e"),
  1322 => (x"6e",x"51",x"66",x"d4"),
  1323 => (x"dc",x"81",x"ca",x"49"),
  1324 => (x"66",x"d0",x"51",x"66"),
  1325 => (x"d4",x"80",x"c1",x"48"),
  1326 => (x"66",x"c8",x"58",x"a6"),
  1327 => (x"a8",x"66",x"cc",x"48"),
  1328 => (x"87",x"cb",x"c0",x"04"),
  1329 => (x"c1",x"48",x"66",x"c8"),
  1330 => (x"58",x"a6",x"cc",x"80"),
  1331 => (x"cc",x"87",x"d9",x"c5"),
  1332 => (x"88",x"c1",x"48",x"66"),
  1333 => (x"c5",x"58",x"a6",x"d0"),
  1334 => (x"dd",x"ff",x"87",x"ce"),
  1335 => (x"e8",x"c0",x"87",x"d1"),
  1336 => (x"dd",x"ff",x"58",x"a6"),
  1337 => (x"e0",x"c0",x"87",x"c9"),
  1338 => (x"ec",x"c0",x"58",x"a6"),
  1339 => (x"ca",x"c0",x"05",x"a8"),
  1340 => (x"48",x"a6",x"dc",x"87"),
  1341 => (x"78",x"66",x"e4",x"c0"),
  1342 => (x"ff",x"87",x"c4",x"c0"),
  1343 => (x"c8",x"87",x"fd",x"d9"),
  1344 => (x"91",x"cb",x"49",x"66"),
  1345 => (x"48",x"66",x"fc",x"c0"),
  1346 => (x"7e",x"70",x"80",x"71"),
  1347 => (x"6e",x"82",x"c8",x"4a"),
  1348 => (x"c0",x"81",x"ca",x"49"),
  1349 => (x"dc",x"51",x"66",x"e4"),
  1350 => (x"81",x"c1",x"49",x"66"),
  1351 => (x"89",x"66",x"e4",x"c0"),
  1352 => (x"30",x"71",x"48",x"c1"),
  1353 => (x"89",x"c1",x"49",x"70"),
  1354 => (x"c2",x"7a",x"97",x"71"),
  1355 => (x"49",x"bf",x"c8",x"de"),
  1356 => (x"29",x"66",x"e4",x"c0"),
  1357 => (x"48",x"4a",x"6a",x"97"),
  1358 => (x"ec",x"c0",x"98",x"71"),
  1359 => (x"49",x"6e",x"58",x"a6"),
  1360 => (x"4d",x"69",x"81",x"c4"),
  1361 => (x"c4",x"48",x"66",x"d8"),
  1362 => (x"c0",x"02",x"a8",x"66"),
  1363 => (x"a6",x"c4",x"87",x"c8"),
  1364 => (x"c0",x"78",x"c0",x"48"),
  1365 => (x"a6",x"c4",x"87",x"c5"),
  1366 => (x"c4",x"78",x"c1",x"48"),
  1367 => (x"e0",x"c0",x"1e",x"66"),
  1368 => (x"ff",x"49",x"75",x"1e"),
  1369 => (x"c8",x"87",x"d9",x"d9"),
  1370 => (x"c0",x"4c",x"70",x"86"),
  1371 => (x"c1",x"06",x"ac",x"b7"),
  1372 => (x"85",x"74",x"87",x"d4"),
  1373 => (x"74",x"49",x"e0",x"c0"),
  1374 => (x"c1",x"4b",x"75",x"89"),
  1375 => (x"71",x"4a",x"c3",x"da"),
  1376 => (x"87",x"e3",x"ec",x"fe"),
  1377 => (x"e0",x"c0",x"85",x"c2"),
  1378 => (x"80",x"c1",x"48",x"66"),
  1379 => (x"58",x"a6",x"e4",x"c0"),
  1380 => (x"49",x"66",x"e8",x"c0"),
  1381 => (x"a9",x"70",x"81",x"c1"),
  1382 => (x"87",x"c8",x"c0",x"02"),
  1383 => (x"c0",x"48",x"a6",x"c4"),
  1384 => (x"87",x"c5",x"c0",x"78"),
  1385 => (x"c1",x"48",x"a6",x"c4"),
  1386 => (x"1e",x"66",x"c4",x"78"),
  1387 => (x"c0",x"49",x"a4",x"c2"),
  1388 => (x"88",x"71",x"48",x"e0"),
  1389 => (x"75",x"1e",x"49",x"70"),
  1390 => (x"c3",x"d8",x"ff",x"49"),
  1391 => (x"c0",x"86",x"c8",x"87"),
  1392 => (x"ff",x"01",x"a8",x"b7"),
  1393 => (x"e0",x"c0",x"87",x"c0"),
  1394 => (x"d1",x"c0",x"02",x"66"),
  1395 => (x"c9",x"49",x"6e",x"87"),
  1396 => (x"66",x"e0",x"c0",x"81"),
  1397 => (x"c1",x"48",x"6e",x"51"),
  1398 => (x"c0",x"78",x"dd",x"c4"),
  1399 => (x"49",x"6e",x"87",x"cc"),
  1400 => (x"51",x"c2",x"81",x"c9"),
  1401 => (x"c6",x"c1",x"48",x"6e"),
  1402 => (x"66",x"c8",x"78",x"c9"),
  1403 => (x"a8",x"66",x"cc",x"48"),
  1404 => (x"87",x"cb",x"c0",x"04"),
  1405 => (x"c1",x"48",x"66",x"c8"),
  1406 => (x"58",x"a6",x"cc",x"80"),
  1407 => (x"cc",x"87",x"e9",x"c0"),
  1408 => (x"88",x"c1",x"48",x"66"),
  1409 => (x"c0",x"58",x"a6",x"d0"),
  1410 => (x"d6",x"ff",x"87",x"de"),
  1411 => (x"4c",x"70",x"87",x"de"),
  1412 => (x"c1",x"87",x"d5",x"c0"),
  1413 => (x"c0",x"05",x"ac",x"c6"),
  1414 => (x"66",x"d0",x"87",x"c8"),
  1415 => (x"d4",x"80",x"c1",x"48"),
  1416 => (x"d6",x"ff",x"58",x"a6"),
  1417 => (x"4c",x"70",x"87",x"c6"),
  1418 => (x"c1",x"48",x"66",x"d4"),
  1419 => (x"58",x"a6",x"d8",x"80"),
  1420 => (x"c0",x"02",x"9c",x"74"),
  1421 => (x"66",x"c8",x"87",x"cb"),
  1422 => (x"66",x"c4",x"c1",x"48"),
  1423 => (x"fe",x"f2",x"04",x"a8"),
  1424 => (x"de",x"d5",x"ff",x"87"),
  1425 => (x"48",x"66",x"c8",x"87"),
  1426 => (x"c0",x"03",x"a8",x"c7"),
  1427 => (x"da",x"c2",x"87",x"e5"),
  1428 => (x"78",x"c0",x"48",x"dc"),
  1429 => (x"cb",x"49",x"66",x"c8"),
  1430 => (x"66",x"fc",x"c0",x"91"),
  1431 => (x"4a",x"a1",x"c4",x"81"),
  1432 => (x"52",x"c0",x"4a",x"6a"),
  1433 => (x"48",x"66",x"c8",x"79"),
  1434 => (x"a6",x"cc",x"80",x"c1"),
  1435 => (x"04",x"a8",x"c7",x"58"),
  1436 => (x"ff",x"87",x"db",x"ff"),
  1437 => (x"df",x"ff",x"8e",x"d4"),
  1438 => (x"6f",x"4c",x"87",x"c9"),
  1439 => (x"2a",x"20",x"64",x"61"),
  1440 => (x"3a",x"00",x"20",x"2e"),
  1441 => (x"73",x"1e",x"00",x"20"),
  1442 => (x"9b",x"4b",x"71",x"1e"),
  1443 => (x"c2",x"87",x"c6",x"02"),
  1444 => (x"c0",x"48",x"d8",x"da"),
  1445 => (x"c2",x"1e",x"c7",x"78"),
  1446 => (x"1e",x"bf",x"d8",x"da"),
  1447 => (x"1e",x"ef",x"dd",x"c1"),
  1448 => (x"bf",x"c0",x"da",x"c2"),
  1449 => (x"87",x"c1",x"ee",x"49"),
  1450 => (x"da",x"c2",x"86",x"cc"),
  1451 => (x"e2",x"49",x"bf",x"c0"),
  1452 => (x"9b",x"73",x"87",x"f9"),
  1453 => (x"c1",x"87",x"c8",x"02"),
  1454 => (x"c0",x"49",x"ef",x"dd"),
  1455 => (x"ff",x"87",x"e0",x"e2"),
  1456 => (x"1e",x"87",x"c4",x"de"),
  1457 => (x"48",x"db",x"dd",x"c1"),
  1458 => (x"df",x"c1",x"50",x"c0"),
  1459 => (x"ff",x"49",x"bf",x"d2"),
  1460 => (x"c0",x"87",x"e4",x"d8"),
  1461 => (x"1e",x"4f",x"26",x"48"),
  1462 => (x"c1",x"87",x"db",x"c7"),
  1463 => (x"87",x"e6",x"fe",x"49"),
  1464 => (x"87",x"cc",x"ef",x"fe"),
  1465 => (x"cd",x"02",x"98",x"70"),
  1466 => (x"e6",x"f6",x"fe",x"87"),
  1467 => (x"02",x"98",x"70",x"87"),
  1468 => (x"4a",x"c1",x"87",x"c4"),
  1469 => (x"4a",x"c0",x"87",x"c2"),
  1470 => (x"ce",x"05",x"9a",x"72"),
  1471 => (x"c1",x"1e",x"c0",x"87"),
  1472 => (x"c0",x"49",x"f2",x"dc"),
  1473 => (x"c4",x"87",x"db",x"ee"),
  1474 => (x"c2",x"87",x"fe",x"86"),
  1475 => (x"c0",x"48",x"d8",x"da"),
  1476 => (x"c0",x"da",x"c2",x"78"),
  1477 => (x"1e",x"78",x"c0",x"48"),
  1478 => (x"49",x"fd",x"dc",x"c1"),
  1479 => (x"87",x"c2",x"ee",x"c0"),
  1480 => (x"de",x"fe",x"1e",x"c0"),
  1481 => (x"c0",x"49",x"70",x"87"),
  1482 => (x"c3",x"87",x"f7",x"ed"),
  1483 => (x"8e",x"f8",x"87",x"c7"),
  1484 => (x"44",x"53",x"4f",x"26"),
  1485 => (x"69",x"61",x"66",x"20"),
  1486 => (x"2e",x"64",x"65",x"6c"),
  1487 => (x"6f",x"6f",x"42",x"00"),
  1488 => (x"67",x"6e",x"69",x"74"),
  1489 => (x"00",x"2e",x"2e",x"2e"),
  1490 => (x"cf",x"e2",x"c0",x"1e"),
  1491 => (x"26",x"87",x"fa",x"87"),
  1492 => (x"c2",x"fe",x"1e",x"4f"),
  1493 => (x"c0",x"87",x"f1",x"87"),
  1494 => (x"00",x"4f",x"26",x"48"),
  1495 => (x"00",x"00",x"01",x"00"),
  1496 => (x"45",x"20",x"80",x"00"),
  1497 => (x"00",x"74",x"69",x"78"),
  1498 => (x"61",x"42",x"20",x"80"),
  1499 => (x"99",x"00",x"6b",x"63"),
  1500 => (x"ac",x"00",x"00",x"0e"),
  1501 => (x"00",x"00",x"00",x"26"),
  1502 => (x"0e",x"99",x"00",x"00"),
  1503 => (x"26",x"ca",x"00",x"00"),
  1504 => (x"00",x"00",x"00",x"00"),
  1505 => (x"00",x"0e",x"99",x"00"),
  1506 => (x"00",x"26",x"e8",x"00"),
  1507 => (x"00",x"00",x"00",x"00"),
  1508 => (x"00",x"00",x"0e",x"99"),
  1509 => (x"00",x"00",x"27",x"06"),
  1510 => (x"99",x"00",x"00",x"00"),
  1511 => (x"24",x"00",x"00",x"0e"),
  1512 => (x"00",x"00",x"00",x"27"),
  1513 => (x"0e",x"99",x"00",x"00"),
  1514 => (x"27",x"42",x"00",x"00"),
  1515 => (x"00",x"00",x"00",x"00"),
  1516 => (x"00",x"0e",x"99",x"00"),
  1517 => (x"00",x"27",x"60",x"00"),
  1518 => (x"00",x"00",x"00",x"00"),
  1519 => (x"00",x"00",x"0f",x"4c"),
  1520 => (x"00",x"00",x"00",x"00"),
  1521 => (x"9a",x"00",x"00",x"00"),
  1522 => (x"00",x"00",x"00",x"11"),
  1523 => (x"00",x"00",x"00",x"00"),
  1524 => (x"17",x"d6",x"00",x"00"),
  1525 => (x"4f",x"42",x"00",x"00"),
  1526 => (x"20",x"20",x"54",x"4f"),
  1527 => (x"4f",x"52",x"20",x"20"),
  1528 => (x"fe",x"1e",x"00",x"4d"),
  1529 => (x"78",x"c0",x"48",x"f0"),
  1530 => (x"09",x"79",x"09",x"cd"),
  1531 => (x"fe",x"1e",x"4f",x"26"),
  1532 => (x"26",x"48",x"bf",x"f0"),
  1533 => (x"f0",x"fe",x"1e",x"4f"),
  1534 => (x"26",x"78",x"c1",x"48"),
  1535 => (x"f0",x"fe",x"1e",x"4f"),
  1536 => (x"26",x"78",x"c0",x"48"),
  1537 => (x"4a",x"71",x"1e",x"4f"),
  1538 => (x"26",x"52",x"52",x"c0"),
  1539 => (x"5b",x"5e",x"0e",x"4f"),
  1540 => (x"f4",x"0e",x"5d",x"5c"),
  1541 => (x"97",x"4d",x"71",x"86"),
  1542 => (x"a5",x"c1",x"7e",x"6d"),
  1543 => (x"48",x"6c",x"97",x"4c"),
  1544 => (x"6e",x"58",x"a6",x"c8"),
  1545 => (x"a8",x"66",x"c4",x"48"),
  1546 => (x"ff",x"87",x"c5",x"05"),
  1547 => (x"87",x"e6",x"c0",x"48"),
  1548 => (x"c2",x"87",x"ca",x"ff"),
  1549 => (x"6c",x"97",x"49",x"a5"),
  1550 => (x"4b",x"a3",x"71",x"4b"),
  1551 => (x"97",x"4b",x"6b",x"97"),
  1552 => (x"48",x"6e",x"7e",x"6c"),
  1553 => (x"a6",x"c8",x"80",x"c1"),
  1554 => (x"cc",x"98",x"c7",x"58"),
  1555 => (x"97",x"70",x"58",x"a6"),
  1556 => (x"87",x"e1",x"fe",x"7c"),
  1557 => (x"8e",x"f4",x"48",x"73"),
  1558 => (x"4c",x"26",x"4d",x"26"),
  1559 => (x"4f",x"26",x"4b",x"26"),
  1560 => (x"5c",x"5b",x"5e",x"0e"),
  1561 => (x"71",x"86",x"f4",x"0e"),
  1562 => (x"4a",x"66",x"d8",x"4c"),
  1563 => (x"c2",x"9a",x"ff",x"c3"),
  1564 => (x"6c",x"97",x"4b",x"a4"),
  1565 => (x"49",x"a1",x"73",x"49"),
  1566 => (x"6c",x"97",x"51",x"72"),
  1567 => (x"c1",x"48",x"6e",x"7e"),
  1568 => (x"58",x"a6",x"c8",x"80"),
  1569 => (x"a6",x"cc",x"98",x"c7"),
  1570 => (x"f4",x"54",x"70",x"58"),
  1571 => (x"87",x"ca",x"ff",x"8e"),
  1572 => (x"e8",x"fd",x"1e",x"1e"),
  1573 => (x"4a",x"bf",x"e0",x"87"),
  1574 => (x"c0",x"e0",x"c0",x"49"),
  1575 => (x"87",x"cb",x"02",x"99"),
  1576 => (x"dd",x"c2",x"1e",x"72"),
  1577 => (x"f7",x"fe",x"49",x"fe"),
  1578 => (x"fd",x"86",x"c4",x"87"),
  1579 => (x"7e",x"70",x"87",x"c0"),
  1580 => (x"26",x"87",x"c2",x"fd"),
  1581 => (x"c2",x"1e",x"4f",x"26"),
  1582 => (x"fd",x"49",x"fe",x"dd"),
  1583 => (x"e2",x"c1",x"87",x"c7"),
  1584 => (x"dd",x"fc",x"49",x"d0"),
  1585 => (x"87",x"ee",x"c3",x"87"),
  1586 => (x"5e",x"0e",x"4f",x"26"),
  1587 => (x"0e",x"5d",x"5c",x"5b"),
  1588 => (x"dd",x"c2",x"4d",x"71"),
  1589 => (x"f4",x"fc",x"49",x"fe"),
  1590 => (x"c0",x"4b",x"70",x"87"),
  1591 => (x"c3",x"04",x"ab",x"b7"),
  1592 => (x"f0",x"c3",x"87",x"c2"),
  1593 => (x"87",x"c9",x"05",x"ab"),
  1594 => (x"48",x"ee",x"e6",x"c1"),
  1595 => (x"e3",x"c2",x"78",x"c1"),
  1596 => (x"ab",x"e0",x"c3",x"87"),
  1597 => (x"c1",x"87",x"c9",x"05"),
  1598 => (x"c1",x"48",x"f2",x"e6"),
  1599 => (x"87",x"d4",x"c2",x"78"),
  1600 => (x"bf",x"f2",x"e6",x"c1"),
  1601 => (x"c2",x"87",x"c6",x"02"),
  1602 => (x"c2",x"4c",x"a3",x"c0"),
  1603 => (x"c1",x"4c",x"73",x"87"),
  1604 => (x"02",x"bf",x"ee",x"e6"),
  1605 => (x"74",x"87",x"e0",x"c0"),
  1606 => (x"29",x"b7",x"c4",x"49"),
  1607 => (x"c5",x"e8",x"c1",x"91"),
  1608 => (x"cf",x"4a",x"74",x"81"),
  1609 => (x"c1",x"92",x"c2",x"9a"),
  1610 => (x"70",x"30",x"72",x"48"),
  1611 => (x"72",x"ba",x"ff",x"4a"),
  1612 => (x"70",x"98",x"69",x"48"),
  1613 => (x"74",x"87",x"db",x"79"),
  1614 => (x"29",x"b7",x"c4",x"49"),
  1615 => (x"c5",x"e8",x"c1",x"91"),
  1616 => (x"cf",x"4a",x"74",x"81"),
  1617 => (x"c3",x"92",x"c2",x"9a"),
  1618 => (x"70",x"30",x"72",x"48"),
  1619 => (x"b0",x"69",x"48",x"4a"),
  1620 => (x"9d",x"75",x"79",x"70"),
  1621 => (x"87",x"f0",x"c0",x"05"),
  1622 => (x"c8",x"48",x"d0",x"ff"),
  1623 => (x"d4",x"ff",x"78",x"e1"),
  1624 => (x"c1",x"78",x"c5",x"48"),
  1625 => (x"02",x"bf",x"f2",x"e6"),
  1626 => (x"e0",x"c3",x"87",x"c3"),
  1627 => (x"ee",x"e6",x"c1",x"78"),
  1628 => (x"87",x"c6",x"02",x"bf"),
  1629 => (x"c3",x"48",x"d4",x"ff"),
  1630 => (x"d4",x"ff",x"78",x"f0"),
  1631 => (x"ff",x"0b",x"7b",x"0b"),
  1632 => (x"e1",x"c8",x"48",x"d0"),
  1633 => (x"78",x"e0",x"c0",x"78"),
  1634 => (x"48",x"f2",x"e6",x"c1"),
  1635 => (x"e6",x"c1",x"78",x"c0"),
  1636 => (x"78",x"c0",x"48",x"ee"),
  1637 => (x"49",x"fe",x"dd",x"c2"),
  1638 => (x"70",x"87",x"f2",x"f9"),
  1639 => (x"ab",x"b7",x"c0",x"4b"),
  1640 => (x"87",x"fe",x"fc",x"03"),
  1641 => (x"4d",x"26",x"48",x"c0"),
  1642 => (x"4b",x"26",x"4c",x"26"),
  1643 => (x"00",x"00",x"4f",x"26"),
  1644 => (x"00",x"00",x"00",x"00"),
  1645 => (x"c0",x"1e",x"00",x"00"),
  1646 => (x"c4",x"49",x"72",x"4a"),
  1647 => (x"c5",x"e8",x"c1",x"91"),
  1648 => (x"c1",x"79",x"c0",x"81"),
  1649 => (x"aa",x"b7",x"d0",x"82"),
  1650 => (x"26",x"87",x"ee",x"04"),
  1651 => (x"5b",x"5e",x"0e",x"4f"),
  1652 => (x"71",x"0e",x"5d",x"5c"),
  1653 => (x"87",x"e5",x"f8",x"4d"),
  1654 => (x"b7",x"c4",x"4a",x"75"),
  1655 => (x"e8",x"c1",x"92",x"2a"),
  1656 => (x"4c",x"75",x"82",x"c5"),
  1657 => (x"94",x"c2",x"9c",x"cf"),
  1658 => (x"74",x"4b",x"49",x"6a"),
  1659 => (x"c2",x"9b",x"c3",x"2b"),
  1660 => (x"70",x"30",x"74",x"48"),
  1661 => (x"74",x"bc",x"ff",x"4c"),
  1662 => (x"70",x"98",x"71",x"48"),
  1663 => (x"87",x"f5",x"f7",x"7a"),
  1664 => (x"e1",x"fe",x"48",x"73"),
  1665 => (x"00",x"00",x"00",x"87"),
  1666 => (x"00",x"00",x"00",x"00"),
  1667 => (x"00",x"00",x"00",x"00"),
  1668 => (x"00",x"00",x"00",x"00"),
  1669 => (x"00",x"00",x"00",x"00"),
  1670 => (x"00",x"00",x"00",x"00"),
  1671 => (x"00",x"00",x"00",x"00"),
  1672 => (x"00",x"00",x"00",x"00"),
  1673 => (x"00",x"00",x"00",x"00"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"d0",x"ff",x"1e",x"00"),
  1682 => (x"78",x"e1",x"c8",x"48"),
  1683 => (x"d4",x"ff",x"48",x"71"),
  1684 => (x"66",x"c4",x"78",x"08"),
  1685 => (x"08",x"d4",x"ff",x"48"),
  1686 => (x"1e",x"4f",x"26",x"78"),
  1687 => (x"66",x"c4",x"4a",x"71"),
  1688 => (x"49",x"72",x"1e",x"49"),
  1689 => (x"ff",x"87",x"de",x"ff"),
  1690 => (x"e0",x"c0",x"48",x"d0"),
  1691 => (x"4f",x"26",x"26",x"78"),
  1692 => (x"71",x"1e",x"73",x"1e"),
  1693 => (x"49",x"66",x"c8",x"4b"),
  1694 => (x"c1",x"4a",x"73",x"1e"),
  1695 => (x"ff",x"49",x"a2",x"e0"),
  1696 => (x"c4",x"26",x"87",x"d9"),
  1697 => (x"26",x"4d",x"26",x"87"),
  1698 => (x"26",x"4b",x"26",x"4c"),
  1699 => (x"d4",x"ff",x"1e",x"4f"),
  1700 => (x"7a",x"ff",x"c3",x"4a"),
  1701 => (x"c0",x"48",x"d0",x"ff"),
  1702 => (x"7a",x"de",x"78",x"e1"),
  1703 => (x"bf",x"c8",x"de",x"c2"),
  1704 => (x"c8",x"48",x"49",x"7a"),
  1705 => (x"71",x"7a",x"70",x"28"),
  1706 => (x"70",x"28",x"d0",x"48"),
  1707 => (x"d8",x"48",x"71",x"7a"),
  1708 => (x"ff",x"7a",x"70",x"28"),
  1709 => (x"e0",x"c0",x"48",x"d0"),
  1710 => (x"1e",x"4f",x"26",x"78"),
  1711 => (x"c8",x"48",x"d0",x"ff"),
  1712 => (x"48",x"71",x"78",x"c9"),
  1713 => (x"78",x"08",x"d4",x"ff"),
  1714 => (x"71",x"1e",x"4f",x"26"),
  1715 => (x"87",x"eb",x"49",x"4a"),
  1716 => (x"c8",x"48",x"d0",x"ff"),
  1717 => (x"1e",x"4f",x"26",x"78"),
  1718 => (x"4b",x"71",x"1e",x"73"),
  1719 => (x"bf",x"d8",x"de",x"c2"),
  1720 => (x"c2",x"87",x"c3",x"02"),
  1721 => (x"d0",x"ff",x"87",x"eb"),
  1722 => (x"78",x"c9",x"c8",x"48"),
  1723 => (x"e0",x"c0",x"48",x"73"),
  1724 => (x"08",x"d4",x"ff",x"b0"),
  1725 => (x"cc",x"de",x"c2",x"78"),
  1726 => (x"c8",x"78",x"c0",x"48"),
  1727 => (x"87",x"c5",x"02",x"66"),
  1728 => (x"c2",x"49",x"ff",x"c3"),
  1729 => (x"c2",x"49",x"c0",x"87"),
  1730 => (x"cc",x"59",x"d4",x"de"),
  1731 => (x"87",x"c6",x"02",x"66"),
  1732 => (x"4a",x"d5",x"d5",x"c5"),
  1733 => (x"ff",x"cf",x"87",x"c4"),
  1734 => (x"de",x"c2",x"4a",x"ff"),
  1735 => (x"de",x"c2",x"5a",x"d8"),
  1736 => (x"78",x"c1",x"48",x"d8"),
  1737 => (x"4d",x"26",x"87",x"c4"),
  1738 => (x"4b",x"26",x"4c",x"26"),
  1739 => (x"5e",x"0e",x"4f",x"26"),
  1740 => (x"0e",x"5d",x"5c",x"5b"),
  1741 => (x"de",x"c2",x"4a",x"71"),
  1742 => (x"72",x"4c",x"bf",x"d4"),
  1743 => (x"87",x"cb",x"02",x"9a"),
  1744 => (x"c1",x"91",x"c8",x"49"),
  1745 => (x"71",x"4b",x"cd",x"eb"),
  1746 => (x"c1",x"87",x"c4",x"83"),
  1747 => (x"c0",x"4b",x"cd",x"ef"),
  1748 => (x"74",x"49",x"13",x"4d"),
  1749 => (x"d0",x"de",x"c2",x"99"),
  1750 => (x"b8",x"71",x"48",x"bf"),
  1751 => (x"78",x"08",x"d4",x"ff"),
  1752 => (x"85",x"2c",x"b7",x"c1"),
  1753 => (x"04",x"ad",x"b7",x"c8"),
  1754 => (x"de",x"c2",x"87",x"e7"),
  1755 => (x"c8",x"48",x"bf",x"cc"),
  1756 => (x"d0",x"de",x"c2",x"80"),
  1757 => (x"87",x"ee",x"fe",x"58"),
  1758 => (x"71",x"1e",x"73",x"1e"),
  1759 => (x"9a",x"4a",x"13",x"4b"),
  1760 => (x"72",x"87",x"cb",x"02"),
  1761 => (x"87",x"e6",x"fe",x"49"),
  1762 => (x"05",x"9a",x"4a",x"13"),
  1763 => (x"d9",x"fe",x"87",x"f5"),
  1764 => (x"de",x"c2",x"1e",x"87"),
  1765 => (x"c2",x"49",x"bf",x"cc"),
  1766 => (x"c1",x"48",x"cc",x"de"),
  1767 => (x"c0",x"c4",x"78",x"a1"),
  1768 => (x"db",x"03",x"a9",x"b7"),
  1769 => (x"48",x"d4",x"ff",x"87"),
  1770 => (x"bf",x"d0",x"de",x"c2"),
  1771 => (x"cc",x"de",x"c2",x"78"),
  1772 => (x"de",x"c2",x"49",x"bf"),
  1773 => (x"a1",x"c1",x"48",x"cc"),
  1774 => (x"b7",x"c0",x"c4",x"78"),
  1775 => (x"87",x"e5",x"04",x"a9"),
  1776 => (x"c8",x"48",x"d0",x"ff"),
  1777 => (x"d8",x"de",x"c2",x"78"),
  1778 => (x"26",x"78",x"c0",x"48"),
  1779 => (x"00",x"00",x"00",x"4f"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"5f",x"5f"),
  1783 => (x"03",x"03",x"00",x"00"),
  1784 => (x"00",x"03",x"03",x"00"),
  1785 => (x"7f",x"7f",x"14",x"00"),
  1786 => (x"14",x"7f",x"7f",x"14"),
  1787 => (x"2e",x"24",x"00",x"00"),
  1788 => (x"12",x"3a",x"6b",x"6b"),
  1789 => (x"36",x"6a",x"4c",x"00"),
  1790 => (x"32",x"56",x"6c",x"18"),
  1791 => (x"4f",x"7e",x"30",x"00"),
  1792 => (x"68",x"3a",x"77",x"59"),
  1793 => (x"04",x"00",x"00",x"40"),
  1794 => (x"00",x"00",x"03",x"07"),
  1795 => (x"1c",x"00",x"00",x"00"),
  1796 => (x"00",x"41",x"63",x"3e"),
  1797 => (x"41",x"00",x"00",x"00"),
  1798 => (x"00",x"1c",x"3e",x"63"),
  1799 => (x"3e",x"2a",x"08",x"00"),
  1800 => (x"2a",x"3e",x"1c",x"1c"),
  1801 => (x"08",x"08",x"00",x"08"),
  1802 => (x"08",x"08",x"3e",x"3e"),
  1803 => (x"80",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"60",x"e0"),
  1805 => (x"08",x"08",x"00",x"00"),
  1806 => (x"08",x"08",x"08",x"08"),
  1807 => (x"00",x"00",x"00",x"00"),
  1808 => (x"00",x"00",x"60",x"60"),
  1809 => (x"30",x"60",x"40",x"00"),
  1810 => (x"03",x"06",x"0c",x"18"),
  1811 => (x"7f",x"3e",x"00",x"01"),
  1812 => (x"3e",x"7f",x"4d",x"59"),
  1813 => (x"06",x"04",x"00",x"00"),
  1814 => (x"00",x"00",x"7f",x"7f"),
  1815 => (x"63",x"42",x"00",x"00"),
  1816 => (x"46",x"4f",x"59",x"71"),
  1817 => (x"63",x"22",x"00",x"00"),
  1818 => (x"36",x"7f",x"49",x"49"),
  1819 => (x"16",x"1c",x"18",x"00"),
  1820 => (x"10",x"7f",x"7f",x"13"),
  1821 => (x"67",x"27",x"00",x"00"),
  1822 => (x"39",x"7d",x"45",x"45"),
  1823 => (x"7e",x"3c",x"00",x"00"),
  1824 => (x"30",x"79",x"49",x"4b"),
  1825 => (x"01",x"01",x"00",x"00"),
  1826 => (x"07",x"0f",x"79",x"71"),
  1827 => (x"7f",x"36",x"00",x"00"),
  1828 => (x"36",x"7f",x"49",x"49"),
  1829 => (x"4f",x"06",x"00",x"00"),
  1830 => (x"1e",x"3f",x"69",x"49"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"66",x"66"),
  1833 => (x"80",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"66",x"e6"),
  1835 => (x"08",x"08",x"00",x"00"),
  1836 => (x"22",x"22",x"14",x"14"),
  1837 => (x"14",x"14",x"00",x"00"),
  1838 => (x"14",x"14",x"14",x"14"),
  1839 => (x"22",x"22",x"00",x"00"),
  1840 => (x"08",x"08",x"14",x"14"),
  1841 => (x"03",x"02",x"00",x"00"),
  1842 => (x"06",x"0f",x"59",x"51"),
  1843 => (x"41",x"7f",x"3e",x"00"),
  1844 => (x"1e",x"1f",x"55",x"5d"),
  1845 => (x"7f",x"7e",x"00",x"00"),
  1846 => (x"7e",x"7f",x"09",x"09"),
  1847 => (x"7f",x"7f",x"00",x"00"),
  1848 => (x"36",x"7f",x"49",x"49"),
  1849 => (x"3e",x"1c",x"00",x"00"),
  1850 => (x"41",x"41",x"41",x"63"),
  1851 => (x"7f",x"7f",x"00",x"00"),
  1852 => (x"1c",x"3e",x"63",x"41"),
  1853 => (x"7f",x"7f",x"00",x"00"),
  1854 => (x"41",x"41",x"49",x"49"),
  1855 => (x"7f",x"7f",x"00",x"00"),
  1856 => (x"01",x"01",x"09",x"09"),
  1857 => (x"7f",x"3e",x"00",x"00"),
  1858 => (x"7a",x"7b",x"49",x"41"),
  1859 => (x"7f",x"7f",x"00",x"00"),
  1860 => (x"7f",x"7f",x"08",x"08"),
  1861 => (x"41",x"00",x"00",x"00"),
  1862 => (x"00",x"41",x"7f",x"7f"),
  1863 => (x"60",x"20",x"00",x"00"),
  1864 => (x"3f",x"7f",x"40",x"40"),
  1865 => (x"08",x"7f",x"7f",x"00"),
  1866 => (x"41",x"63",x"36",x"1c"),
  1867 => (x"7f",x"7f",x"00",x"00"),
  1868 => (x"40",x"40",x"40",x"40"),
  1869 => (x"06",x"7f",x"7f",x"00"),
  1870 => (x"7f",x"7f",x"06",x"0c"),
  1871 => (x"06",x"7f",x"7f",x"00"),
  1872 => (x"7f",x"7f",x"18",x"0c"),
  1873 => (x"7f",x"3e",x"00",x"00"),
  1874 => (x"3e",x"7f",x"41",x"41"),
  1875 => (x"7f",x"7f",x"00",x"00"),
  1876 => (x"06",x"0f",x"09",x"09"),
  1877 => (x"41",x"7f",x"3e",x"00"),
  1878 => (x"40",x"7e",x"7f",x"61"),
  1879 => (x"7f",x"7f",x"00",x"00"),
  1880 => (x"66",x"7f",x"19",x"09"),
  1881 => (x"6f",x"26",x"00",x"00"),
  1882 => (x"32",x"7b",x"59",x"4d"),
  1883 => (x"01",x"01",x"00",x"00"),
  1884 => (x"01",x"01",x"7f",x"7f"),
  1885 => (x"7f",x"3f",x"00",x"00"),
  1886 => (x"3f",x"7f",x"40",x"40"),
  1887 => (x"3f",x"0f",x"00",x"00"),
  1888 => (x"0f",x"3f",x"70",x"70"),
  1889 => (x"30",x"7f",x"7f",x"00"),
  1890 => (x"7f",x"7f",x"30",x"18"),
  1891 => (x"36",x"63",x"41",x"00"),
  1892 => (x"63",x"36",x"1c",x"1c"),
  1893 => (x"06",x"03",x"01",x"41"),
  1894 => (x"03",x"06",x"7c",x"7c"),
  1895 => (x"59",x"71",x"61",x"01"),
  1896 => (x"41",x"43",x"47",x"4d"),
  1897 => (x"7f",x"00",x"00",x"00"),
  1898 => (x"00",x"41",x"41",x"7f"),
  1899 => (x"06",x"03",x"01",x"00"),
  1900 => (x"60",x"30",x"18",x"0c"),
  1901 => (x"41",x"00",x"00",x"40"),
  1902 => (x"00",x"7f",x"7f",x"41"),
  1903 => (x"06",x"0c",x"08",x"00"),
  1904 => (x"08",x"0c",x"06",x"03"),
  1905 => (x"80",x"80",x"80",x"00"),
  1906 => (x"80",x"80",x"80",x"80"),
  1907 => (x"00",x"00",x"00",x"00"),
  1908 => (x"00",x"04",x"07",x"03"),
  1909 => (x"74",x"20",x"00",x"00"),
  1910 => (x"78",x"7c",x"54",x"54"),
  1911 => (x"7f",x"7f",x"00",x"00"),
  1912 => (x"38",x"7c",x"44",x"44"),
  1913 => (x"7c",x"38",x"00",x"00"),
  1914 => (x"00",x"44",x"44",x"44"),
  1915 => (x"7c",x"38",x"00",x"00"),
  1916 => (x"7f",x"7f",x"44",x"44"),
  1917 => (x"7c",x"38",x"00",x"00"),
  1918 => (x"18",x"5c",x"54",x"54"),
  1919 => (x"7e",x"04",x"00",x"00"),
  1920 => (x"00",x"05",x"05",x"7f"),
  1921 => (x"bc",x"18",x"00",x"00"),
  1922 => (x"7c",x"fc",x"a4",x"a4"),
  1923 => (x"7f",x"7f",x"00",x"00"),
  1924 => (x"78",x"7c",x"04",x"04"),
  1925 => (x"00",x"00",x"00",x"00"),
  1926 => (x"00",x"40",x"7d",x"3d"),
  1927 => (x"80",x"80",x"00",x"00"),
  1928 => (x"00",x"7d",x"fd",x"80"),
  1929 => (x"7f",x"7f",x"00",x"00"),
  1930 => (x"44",x"6c",x"38",x"10"),
  1931 => (x"00",x"00",x"00",x"00"),
  1932 => (x"00",x"40",x"7f",x"3f"),
  1933 => (x"0c",x"7c",x"7c",x"00"),
  1934 => (x"78",x"7c",x"0c",x"18"),
  1935 => (x"7c",x"7c",x"00",x"00"),
  1936 => (x"78",x"7c",x"04",x"04"),
  1937 => (x"7c",x"38",x"00",x"00"),
  1938 => (x"38",x"7c",x"44",x"44"),
  1939 => (x"fc",x"fc",x"00",x"00"),
  1940 => (x"18",x"3c",x"24",x"24"),
  1941 => (x"3c",x"18",x"00",x"00"),
  1942 => (x"fc",x"fc",x"24",x"24"),
  1943 => (x"7c",x"7c",x"00",x"00"),
  1944 => (x"08",x"0c",x"04",x"04"),
  1945 => (x"5c",x"48",x"00",x"00"),
  1946 => (x"20",x"74",x"54",x"54"),
  1947 => (x"3f",x"04",x"00",x"00"),
  1948 => (x"00",x"44",x"44",x"7f"),
  1949 => (x"7c",x"3c",x"00",x"00"),
  1950 => (x"7c",x"7c",x"40",x"40"),
  1951 => (x"3c",x"1c",x"00",x"00"),
  1952 => (x"1c",x"3c",x"60",x"60"),
  1953 => (x"60",x"7c",x"3c",x"00"),
  1954 => (x"3c",x"7c",x"60",x"30"),
  1955 => (x"38",x"6c",x"44",x"00"),
  1956 => (x"44",x"6c",x"38",x"10"),
  1957 => (x"bc",x"1c",x"00",x"00"),
  1958 => (x"1c",x"3c",x"60",x"e0"),
  1959 => (x"64",x"44",x"00",x"00"),
  1960 => (x"44",x"4c",x"5c",x"74"),
  1961 => (x"08",x"08",x"00",x"00"),
  1962 => (x"41",x"41",x"77",x"3e"),
  1963 => (x"00",x"00",x"00",x"00"),
  1964 => (x"00",x"00",x"7f",x"7f"),
  1965 => (x"41",x"41",x"00",x"00"),
  1966 => (x"08",x"08",x"3e",x"77"),
  1967 => (x"01",x"01",x"02",x"00"),
  1968 => (x"01",x"02",x"02",x"03"),
  1969 => (x"7f",x"7f",x"7f",x"00"),
  1970 => (x"7f",x"7f",x"7f",x"7f"),
  1971 => (x"1c",x"08",x"08",x"00"),
  1972 => (x"7f",x"3e",x"3e",x"1c"),
  1973 => (x"3e",x"7f",x"7f",x"7f"),
  1974 => (x"08",x"1c",x"1c",x"3e"),
  1975 => (x"18",x"10",x"00",x"08"),
  1976 => (x"10",x"18",x"7c",x"7c"),
  1977 => (x"30",x"10",x"00",x"00"),
  1978 => (x"10",x"30",x"7c",x"7c"),
  1979 => (x"60",x"30",x"10",x"00"),
  1980 => (x"06",x"1e",x"78",x"60"),
  1981 => (x"3c",x"66",x"42",x"00"),
  1982 => (x"42",x"66",x"3c",x"18"),
  1983 => (x"6a",x"38",x"78",x"00"),
  1984 => (x"38",x"6c",x"c6",x"c2"),
  1985 => (x"00",x"00",x"60",x"00"),
  1986 => (x"60",x"00",x"00",x"60"),
  1987 => (x"5b",x"5e",x"0e",x"00"),
  1988 => (x"1e",x"0e",x"5d",x"5c"),
  1989 => (x"de",x"c2",x"4c",x"71"),
  1990 => (x"c0",x"4d",x"bf",x"dd"),
  1991 => (x"74",x"1e",x"c0",x"4b"),
  1992 => (x"87",x"c7",x"02",x"ab"),
  1993 => (x"c0",x"48",x"a6",x"c4"),
  1994 => (x"c4",x"87",x"c5",x"78"),
  1995 => (x"78",x"c1",x"48",x"a6"),
  1996 => (x"73",x"1e",x"66",x"c4"),
  1997 => (x"87",x"df",x"ee",x"49"),
  1998 => (x"e0",x"c0",x"86",x"c8"),
  1999 => (x"87",x"ee",x"ef",x"49"),
  2000 => (x"6a",x"4a",x"a5",x"c4"),
  2001 => (x"87",x"f0",x"f0",x"49"),
  2002 => (x"cb",x"87",x"c6",x"f1"),
  2003 => (x"c8",x"83",x"c1",x"85"),
  2004 => (x"ff",x"04",x"ab",x"b7"),
  2005 => (x"26",x"26",x"87",x"c7"),
  2006 => (x"26",x"4c",x"26",x"4d"),
  2007 => (x"1e",x"4f",x"26",x"4b"),
  2008 => (x"de",x"c2",x"4a",x"71"),
  2009 => (x"de",x"c2",x"5a",x"e1"),
  2010 => (x"78",x"c7",x"48",x"e1"),
  2011 => (x"87",x"dd",x"fe",x"49"),
  2012 => (x"73",x"1e",x"4f",x"26"),
  2013 => (x"c0",x"4a",x"71",x"1e"),
  2014 => (x"d3",x"03",x"aa",x"b7"),
  2015 => (x"fb",x"cb",x"c2",x"87"),
  2016 => (x"87",x"c4",x"05",x"bf"),
  2017 => (x"87",x"c2",x"4b",x"c1"),
  2018 => (x"cb",x"c2",x"4b",x"c0"),
  2019 => (x"87",x"c4",x"5b",x"ff"),
  2020 => (x"5a",x"ff",x"cb",x"c2"),
  2021 => (x"bf",x"fb",x"cb",x"c2"),
  2022 => (x"c1",x"9a",x"c1",x"4a"),
  2023 => (x"ec",x"49",x"a2",x"c0"),
  2024 => (x"48",x"fc",x"87",x"e8"),
  2025 => (x"bf",x"fb",x"cb",x"c2"),
  2026 => (x"87",x"ef",x"fe",x"78"),
  2027 => (x"c4",x"4a",x"71",x"1e"),
  2028 => (x"49",x"72",x"1e",x"66"),
  2029 => (x"26",x"87",x"f9",x"ea"),
  2030 => (x"ff",x"1e",x"4f",x"26"),
  2031 => (x"ff",x"c3",x"48",x"d4"),
  2032 => (x"48",x"d0",x"ff",x"78"),
  2033 => (x"ff",x"78",x"e1",x"c0"),
  2034 => (x"78",x"c1",x"48",x"d4"),
  2035 => (x"30",x"c4",x"48",x"71"),
  2036 => (x"78",x"08",x"d4",x"ff"),
  2037 => (x"c0",x"48",x"d0",x"ff"),
  2038 => (x"4f",x"26",x"78",x"e0"),
  2039 => (x"5c",x"5b",x"5e",x"0e"),
  2040 => (x"86",x"f0",x"0e",x"5d"),
  2041 => (x"c0",x"48",x"a6",x"c8"),
  2042 => (x"ec",x"4b",x"4d",x"78"),
  2043 => (x"80",x"fc",x"7e",x"bf"),
  2044 => (x"bf",x"dd",x"de",x"c2"),
  2045 => (x"4c",x"bf",x"e8",x"78"),
  2046 => (x"bf",x"fb",x"cb",x"c2"),
  2047 => (x"87",x"ca",x"e3",x"49"),
  2048 => (x"cb",x"49",x"ee",x"cb"),
  2049 => (x"a6",x"d0",x"87",x"fd"),
  2050 => (x"e6",x"49",x"c7",x"58"),
  2051 => (x"98",x"70",x"87",x"ff"),
  2052 => (x"6e",x"87",x"c8",x"05"),
  2053 => (x"02",x"99",x"c1",x"49"),
  2054 => (x"c1",x"87",x"c3",x"c1"),
  2055 => (x"7e",x"bf",x"ec",x"4b"),
  2056 => (x"bf",x"fb",x"cb",x"c2"),
  2057 => (x"87",x"e2",x"e2",x"49"),
  2058 => (x"cb",x"49",x"66",x"cc"),
  2059 => (x"98",x"70",x"87",x"e1"),
  2060 => (x"c2",x"87",x"d8",x"02"),
  2061 => (x"49",x"bf",x"f3",x"cb"),
  2062 => (x"cb",x"c2",x"b9",x"c1"),
  2063 => (x"fd",x"71",x"59",x"f7"),
  2064 => (x"ee",x"cb",x"87",x"f8"),
  2065 => (x"87",x"fb",x"ca",x"49"),
  2066 => (x"c7",x"58",x"a6",x"d0"),
  2067 => (x"87",x"fd",x"e5",x"49"),
  2068 => (x"ff",x"05",x"98",x"70"),
  2069 => (x"49",x"6e",x"87",x"c5"),
  2070 => (x"fe",x"05",x"99",x"c1"),
  2071 => (x"9b",x"73",x"87",x"fd"),
  2072 => (x"ff",x"87",x"d0",x"02"),
  2073 => (x"87",x"ca",x"fc",x"49"),
  2074 => (x"e5",x"49",x"da",x"c1"),
  2075 => (x"a6",x"c8",x"87",x"df"),
  2076 => (x"c2",x"78",x"c1",x"48"),
  2077 => (x"05",x"bf",x"fb",x"cb"),
  2078 => (x"c3",x"87",x"e9",x"c0"),
  2079 => (x"cc",x"e5",x"49",x"fd"),
  2080 => (x"49",x"fa",x"c3",x"87"),
  2081 => (x"74",x"87",x"c6",x"e5"),
  2082 => (x"99",x"ff",x"c3",x"49"),
  2083 => (x"49",x"c0",x"1e",x"71"),
  2084 => (x"74",x"87",x"d9",x"fc"),
  2085 => (x"29",x"b7",x"c8",x"49"),
  2086 => (x"49",x"c1",x"1e",x"71"),
  2087 => (x"c8",x"87",x"cd",x"fc"),
  2088 => (x"87",x"f9",x"c7",x"86"),
  2089 => (x"ff",x"c3",x"49",x"74"),
  2090 => (x"2c",x"b7",x"c8",x"99"),
  2091 => (x"9c",x"74",x"b4",x"71"),
  2092 => (x"c2",x"87",x"dd",x"02"),
  2093 => (x"49",x"bf",x"f7",x"cb"),
  2094 => (x"70",x"87",x"d4",x"c9"),
  2095 => (x"87",x"c4",x"05",x"98"),
  2096 => (x"87",x"d2",x"4c",x"c0"),
  2097 => (x"c8",x"49",x"e0",x"c2"),
  2098 => (x"cb",x"c2",x"87",x"f9"),
  2099 => (x"87",x"c6",x"58",x"fb"),
  2100 => (x"48",x"f7",x"cb",x"c2"),
  2101 => (x"49",x"74",x"78",x"c0"),
  2102 => (x"ce",x"05",x"99",x"c2"),
  2103 => (x"49",x"eb",x"c3",x"87"),
  2104 => (x"70",x"87",x"ea",x"e3"),
  2105 => (x"02",x"99",x"c2",x"49"),
  2106 => (x"fb",x"87",x"c2",x"c0"),
  2107 => (x"c1",x"49",x"74",x"4d"),
  2108 => (x"87",x"ce",x"05",x"99"),
  2109 => (x"e3",x"49",x"f4",x"c3"),
  2110 => (x"49",x"70",x"87",x"d3"),
  2111 => (x"c0",x"02",x"99",x"c2"),
  2112 => (x"4d",x"fa",x"87",x"c2"),
  2113 => (x"99",x"c8",x"49",x"74"),
  2114 => (x"c3",x"87",x"cd",x"05"),
  2115 => (x"fc",x"e2",x"49",x"f5"),
  2116 => (x"c2",x"49",x"70",x"87"),
  2117 => (x"87",x"d9",x"02",x"99"),
  2118 => (x"bf",x"e1",x"de",x"c2"),
  2119 => (x"87",x"ca",x"c0",x"02"),
  2120 => (x"c2",x"88",x"c1",x"48"),
  2121 => (x"c0",x"58",x"e5",x"de"),
  2122 => (x"4d",x"ff",x"87",x"c2"),
  2123 => (x"c1",x"48",x"a6",x"c8"),
  2124 => (x"c4",x"49",x"74",x"78"),
  2125 => (x"cd",x"c0",x"05",x"99"),
  2126 => (x"49",x"f2",x"c3",x"87"),
  2127 => (x"70",x"87",x"ce",x"e2"),
  2128 => (x"02",x"99",x"c2",x"49"),
  2129 => (x"de",x"c2",x"87",x"df"),
  2130 => (x"48",x"7e",x"bf",x"e1"),
  2131 => (x"03",x"a8",x"b7",x"c7"),
  2132 => (x"6e",x"87",x"cb",x"c0"),
  2133 => (x"c2",x"80",x"c1",x"48"),
  2134 => (x"c0",x"58",x"e5",x"de"),
  2135 => (x"4d",x"fe",x"87",x"c2"),
  2136 => (x"c1",x"48",x"a6",x"c8"),
  2137 => (x"49",x"fd",x"c3",x"78"),
  2138 => (x"70",x"87",x"e2",x"e1"),
  2139 => (x"02",x"99",x"c2",x"49"),
  2140 => (x"c2",x"87",x"d8",x"c0"),
  2141 => (x"02",x"bf",x"e1",x"de"),
  2142 => (x"c2",x"87",x"c9",x"c0"),
  2143 => (x"c0",x"48",x"e1",x"de"),
  2144 => (x"87",x"c2",x"c0",x"78"),
  2145 => (x"a6",x"c8",x"4d",x"fd"),
  2146 => (x"c3",x"78",x"c1",x"48"),
  2147 => (x"fc",x"e0",x"49",x"fa"),
  2148 => (x"c2",x"49",x"70",x"87"),
  2149 => (x"dc",x"c0",x"02",x"99"),
  2150 => (x"e1",x"de",x"c2",x"87"),
  2151 => (x"b7",x"c7",x"48",x"bf"),
  2152 => (x"c9",x"c0",x"03",x"a8"),
  2153 => (x"e1",x"de",x"c2",x"87"),
  2154 => (x"c0",x"78",x"c7",x"48"),
  2155 => (x"4d",x"fc",x"87",x"c2"),
  2156 => (x"c1",x"48",x"a6",x"c8"),
  2157 => (x"ad",x"b7",x"c0",x"78"),
  2158 => (x"87",x"d0",x"c0",x"03"),
  2159 => (x"c1",x"4a",x"66",x"c4"),
  2160 => (x"02",x"6a",x"82",x"d8"),
  2161 => (x"4b",x"87",x"c5",x"c0"),
  2162 => (x"0f",x"73",x"49",x"75"),
  2163 => (x"de",x"c2",x"4b",x"c0"),
  2164 => (x"50",x"c0",x"48",x"dc"),
  2165 => (x"c4",x"49",x"ee",x"cb"),
  2166 => (x"a6",x"d0",x"87",x"e9"),
  2167 => (x"dc",x"de",x"c2",x"58"),
  2168 => (x"c1",x"05",x"bf",x"97"),
  2169 => (x"49",x"74",x"87",x"de"),
  2170 => (x"05",x"99",x"f0",x"c3"),
  2171 => (x"c1",x"87",x"cd",x"c0"),
  2172 => (x"df",x"ff",x"49",x"da"),
  2173 => (x"98",x"70",x"87",x"d7"),
  2174 => (x"87",x"c8",x"c1",x"02"),
  2175 => (x"bf",x"e8",x"4b",x"c1"),
  2176 => (x"ff",x"c3",x"49",x"4c"),
  2177 => (x"2c",x"b7",x"c8",x"99"),
  2178 => (x"cb",x"c2",x"b4",x"71"),
  2179 => (x"ff",x"49",x"bf",x"fb"),
  2180 => (x"cc",x"87",x"f7",x"da"),
  2181 => (x"f6",x"c3",x"49",x"66"),
  2182 => (x"02",x"98",x"70",x"87"),
  2183 => (x"c2",x"87",x"c6",x"c0"),
  2184 => (x"c1",x"48",x"dc",x"de"),
  2185 => (x"dc",x"de",x"c2",x"50"),
  2186 => (x"c0",x"05",x"bf",x"97"),
  2187 => (x"49",x"74",x"87",x"d6"),
  2188 => (x"05",x"99",x"f0",x"c3"),
  2189 => (x"c1",x"87",x"c5",x"ff"),
  2190 => (x"de",x"ff",x"49",x"da"),
  2191 => (x"98",x"70",x"87",x"cf"),
  2192 => (x"87",x"f8",x"fe",x"05"),
  2193 => (x"c0",x"02",x"9b",x"73"),
  2194 => (x"a6",x"cc",x"87",x"e0"),
  2195 => (x"e1",x"de",x"c2",x"48"),
  2196 => (x"66",x"cc",x"78",x"bf"),
  2197 => (x"c4",x"91",x"cb",x"49"),
  2198 => (x"80",x"71",x"48",x"66"),
  2199 => (x"bf",x"6e",x"7e",x"70"),
  2200 => (x"87",x"c6",x"c0",x"02"),
  2201 => (x"49",x"66",x"cc",x"4b"),
  2202 => (x"66",x"c8",x"0f",x"73"),
  2203 => (x"87",x"c8",x"c0",x"02"),
  2204 => (x"bf",x"e1",x"de",x"c2"),
  2205 => (x"87",x"d5",x"f2",x"49"),
  2206 => (x"bf",x"ff",x"cb",x"c2"),
  2207 => (x"87",x"dd",x"c0",x"02"),
  2208 => (x"87",x"cb",x"c2",x"49"),
  2209 => (x"c0",x"02",x"98",x"70"),
  2210 => (x"de",x"c2",x"87",x"d3"),
  2211 => (x"f1",x"49",x"bf",x"e1"),
  2212 => (x"49",x"c0",x"87",x"fb"),
  2213 => (x"c2",x"87",x"db",x"f3"),
  2214 => (x"c0",x"48",x"ff",x"cb"),
  2215 => (x"f2",x"8e",x"f0",x"78"),
  2216 => (x"5e",x"0e",x"87",x"f5"),
  2217 => (x"0e",x"5d",x"5c",x"5b"),
  2218 => (x"c2",x"4c",x"71",x"1e"),
  2219 => (x"49",x"bf",x"dd",x"de"),
  2220 => (x"4d",x"a1",x"cd",x"c1"),
  2221 => (x"69",x"81",x"d1",x"c1"),
  2222 => (x"02",x"9c",x"74",x"7e"),
  2223 => (x"a5",x"c4",x"87",x"cf"),
  2224 => (x"c2",x"7b",x"74",x"4b"),
  2225 => (x"49",x"bf",x"dd",x"de"),
  2226 => (x"6e",x"87",x"d4",x"f2"),
  2227 => (x"05",x"9c",x"74",x"7b"),
  2228 => (x"4b",x"c0",x"87",x"c4"),
  2229 => (x"4b",x"c1",x"87",x"c2"),
  2230 => (x"d5",x"f2",x"49",x"73"),
  2231 => (x"02",x"66",x"d4",x"87"),
  2232 => (x"de",x"49",x"87",x"c7"),
  2233 => (x"c2",x"4a",x"70",x"87"),
  2234 => (x"c2",x"4a",x"c0",x"87"),
  2235 => (x"26",x"5a",x"c3",x"cc"),
  2236 => (x"00",x"87",x"e4",x"f1"),
  2237 => (x"00",x"00",x"00",x"00"),
  2238 => (x"00",x"00",x"00",x"00"),
  2239 => (x"00",x"00",x"00",x"00"),
  2240 => (x"1e",x"00",x"00",x"00"),
  2241 => (x"c8",x"ff",x"4a",x"71"),
  2242 => (x"a1",x"72",x"49",x"bf"),
  2243 => (x"1e",x"4f",x"26",x"48"),
  2244 => (x"89",x"bf",x"c8",x"ff"),
  2245 => (x"c0",x"c0",x"c0",x"fe"),
  2246 => (x"01",x"a9",x"c0",x"c0"),
  2247 => (x"4a",x"c0",x"87",x"c4"),
  2248 => (x"4a",x"c1",x"87",x"c2"),
  2249 => (x"4f",x"26",x"48",x"72"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

