library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0dec287",
    12 => x"86c0c84e",
    13 => x"49f0dec2",
    14 => x"48f0ccc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cbdc",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c348724c",
    72 => x"7c7098ff",
    73 => x"bff0ccc2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"ffc34871",
    79 => x"d07c7098",
    80 => x"29d04966",
    81 => x"ffc34871",
    82 => x"d07c7098",
    83 => x"29c84966",
    84 => x"ffc34871",
    85 => x"d07c7098",
    86 => x"ffc34866",
    87 => x"727c7098",
    88 => x"7129d049",
    89 => x"98ffc348",
    90 => x"4b6c7c70",
    91 => x"4dfff0c9",
    92 => x"05abffc3",
    93 => x"ffc387d0",
    94 => x"c14b6c7c",
    95 => x"87c6028d",
    96 => x"02abffc3",
    97 => x"487387f0",
    98 => x"1e87fffd",
    99 => x"d4ff49c0",
   100 => x"78ffc348",
   101 => x"c8c381c1",
   102 => x"f104a9b7",
   103 => x"1e4f2687",
   104 => x"87e71e73",
   105 => x"4bdff8c4",
   106 => x"ffc01ec0",
   107 => x"49f7c1f0",
   108 => x"c487dffd",
   109 => x"05a8c186",
   110 => x"ff87eac0",
   111 => x"ffc348d4",
   112 => x"c0c0c178",
   113 => x"1ec0c0c0",
   114 => x"c1f0e1c0",
   115 => x"c1fd49e9",
   116 => x"7086c487",
   117 => x"87ca0598",
   118 => x"c348d4ff",
   119 => x"48c178ff",
   120 => x"e6fe87cb",
   121 => x"058bc187",
   122 => x"c087fdfe",
   123 => x"87defc48",
   124 => x"ff1e731e",
   125 => x"ffc348d4",
   126 => x"c04bd378",
   127 => x"f0ffc01e",
   128 => x"fc49c1c1",
   129 => x"86c487cc",
   130 => x"ca059870",
   131 => x"48d4ff87",
   132 => x"c178ffc3",
   133 => x"fd87cb48",
   134 => x"8bc187f1",
   135 => x"87dbff05",
   136 => x"e9fb48c0",
   137 => x"5b5e0e87",
   138 => x"d4ff0e5c",
   139 => x"87dbfd4c",
   140 => x"c01eeac6",
   141 => x"c8c1f0e1",
   142 => x"87d6fb49",
   143 => x"a8c186c4",
   144 => x"fe87c802",
   145 => x"48c087ea",
   146 => x"fa87e2c1",
   147 => x"497087d2",
   148 => x"99ffffcf",
   149 => x"02a9eac6",
   150 => x"d3fe87c8",
   151 => x"c148c087",
   152 => x"ffc387cb",
   153 => x"4bf1c07c",
   154 => x"7087f4fc",
   155 => x"ebc00298",
   156 => x"c01ec087",
   157 => x"fac1f0ff",
   158 => x"87d6fa49",
   159 => x"987086c4",
   160 => x"c387d905",
   161 => x"496c7cff",
   162 => x"7c7cffc3",
   163 => x"c0c17c7c",
   164 => x"87c40299",
   165 => x"87d548c1",
   166 => x"87d148c0",
   167 => x"c405abc2",
   168 => x"c848c087",
   169 => x"058bc187",
   170 => x"c087fdfe",
   171 => x"87dcf948",
   172 => x"c21e731e",
   173 => x"c148f0cc",
   174 => x"ff4bc778",
   175 => x"78c248d0",
   176 => x"ff87c8fb",
   177 => x"78c348d0",
   178 => x"e5c01ec0",
   179 => x"49c0c1d0",
   180 => x"c487fff8",
   181 => x"05a8c186",
   182 => x"c24b87c1",
   183 => x"87c505ab",
   184 => x"f9c048c0",
   185 => x"058bc187",
   186 => x"fc87d0ff",
   187 => x"ccc287f7",
   188 => x"987058f4",
   189 => x"c187cd05",
   190 => x"f0ffc01e",
   191 => x"f849d0c1",
   192 => x"86c487d0",
   193 => x"c348d4ff",
   194 => x"fdc278ff",
   195 => x"f8ccc287",
   196 => x"48d0ff58",
   197 => x"d4ff78c2",
   198 => x"78ffc348",
   199 => x"edf748c1",
   200 => x"5b5e0e87",
   201 => x"710e5d5c",
   202 => x"c54cc04b",
   203 => x"4adfcdee",
   204 => x"c348d4ff",
   205 => x"486878ff",
   206 => x"05a8fec3",
   207 => x"ff87fec0",
   208 => x"9b734dd4",
   209 => x"d087cc02",
   210 => x"49731e66",
   211 => x"c487e8f5",
   212 => x"ff87d686",
   213 => x"d1c448d0",
   214 => x"7dffc378",
   215 => x"c14866d0",
   216 => x"58a6d488",
   217 => x"f0059870",
   218 => x"48d4ff87",
   219 => x"7878ffc3",
   220 => x"c5059b73",
   221 => x"48d0ff87",
   222 => x"4ac178d0",
   223 => x"058ac14c",
   224 => x"7487edfe",
   225 => x"87c2f648",
   226 => x"711e731e",
   227 => x"ff4bc04a",
   228 => x"ffc348d4",
   229 => x"48d0ff78",
   230 => x"ff78c3c4",
   231 => x"ffc348d4",
   232 => x"c01e7278",
   233 => x"d1c1f0ff",
   234 => x"87e6f549",
   235 => x"987086c4",
   236 => x"c887d205",
   237 => x"66cc1ec0",
   238 => x"87e5fd49",
   239 => x"4b7086c4",
   240 => x"c248d0ff",
   241 => x"f5487378",
   242 => x"5e0e87c4",
   243 => x"0e5d5c5b",
   244 => x"ffc01ec0",
   245 => x"49c9c1f0",
   246 => x"d287f7f4",
   247 => x"f8ccc21e",
   248 => x"87fdfc49",
   249 => x"4cc086c8",
   250 => x"b7d284c1",
   251 => x"87f804ac",
   252 => x"97f8ccc2",
   253 => x"c0c349bf",
   254 => x"a9c0c199",
   255 => x"87e7c005",
   256 => x"97ffccc2",
   257 => x"31d049bf",
   258 => x"97c0cdc2",
   259 => x"32c84abf",
   260 => x"cdc2b172",
   261 => x"4abf97c1",
   262 => x"cf4c71b1",
   263 => x"9cffffff",
   264 => x"34ca84c1",
   265 => x"c287e7c1",
   266 => x"bf97c1cd",
   267 => x"c631c149",
   268 => x"c2cdc299",
   269 => x"c74abf97",
   270 => x"b1722ab7",
   271 => x"97fdccc2",
   272 => x"cf4d4abf",
   273 => x"feccc29d",
   274 => x"c34abf97",
   275 => x"c232ca9a",
   276 => x"bf97ffcc",
   277 => x"7333c24b",
   278 => x"c0cdc2b2",
   279 => x"c34bbf97",
   280 => x"b7c69bc0",
   281 => x"c2b2732b",
   282 => x"7148c181",
   283 => x"c1497030",
   284 => x"70307548",
   285 => x"c14c724d",
   286 => x"c8947184",
   287 => x"06adb7c0",
   288 => x"34c187cc",
   289 => x"c0c82db7",
   290 => x"ff01adb7",
   291 => x"487487f4",
   292 => x"0e87f7f1",
   293 => x"5d5c5b5e",
   294 => x"c286f80e",
   295 => x"c048ded5",
   296 => x"d6cdc278",
   297 => x"fb49c01e",
   298 => x"86c487de",
   299 => x"c5059870",
   300 => x"c948c087",
   301 => x"4dc087c0",
   302 => x"edc07ec1",
   303 => x"c249bfeb",
   304 => x"714accce",
   305 => x"e0ee4bc8",
   306 => x"05987087",
   307 => x"7ec087c2",
   308 => x"bfe7edc0",
   309 => x"e8cec249",
   310 => x"4bc8714a",
   311 => x"7087caee",
   312 => x"87c20598",
   313 => x"026e7ec0",
   314 => x"c287fdc0",
   315 => x"4dbfdcd4",
   316 => x"9fd4d5c2",
   317 => x"c5487ebf",
   318 => x"05a8ead6",
   319 => x"d4c287c7",
   320 => x"ce4dbfdc",
   321 => x"ca486e87",
   322 => x"02a8d5e9",
   323 => x"48c087c5",
   324 => x"c287e3c7",
   325 => x"751ed6cd",
   326 => x"87ecf949",
   327 => x"987086c4",
   328 => x"c087c505",
   329 => x"87cec748",
   330 => x"bfe7edc0",
   331 => x"e8cec249",
   332 => x"4bc8714a",
   333 => x"7087f2ec",
   334 => x"87c80598",
   335 => x"48ded5c2",
   336 => x"87da78c1",
   337 => x"bfebedc0",
   338 => x"cccec249",
   339 => x"4bc8714a",
   340 => x"7087d6ec",
   341 => x"c5c00298",
   342 => x"c648c087",
   343 => x"d5c287d8",
   344 => x"49bf97d4",
   345 => x"05a9d5c1",
   346 => x"c287cdc0",
   347 => x"bf97d5d5",
   348 => x"a9eac249",
   349 => x"87c5c002",
   350 => x"f9c548c0",
   351 => x"d6cdc287",
   352 => x"487ebf97",
   353 => x"02a8e9c3",
   354 => x"6e87cec0",
   355 => x"a8ebc348",
   356 => x"87c5c002",
   357 => x"ddc548c0",
   358 => x"e1cdc287",
   359 => x"9949bf97",
   360 => x"87ccc005",
   361 => x"97e2cdc2",
   362 => x"a9c249bf",
   363 => x"87c5c002",
   364 => x"c1c548c0",
   365 => x"e3cdc287",
   366 => x"c248bf97",
   367 => x"7058dad5",
   368 => x"88c1484c",
   369 => x"58ded5c2",
   370 => x"97e4cdc2",
   371 => x"817549bf",
   372 => x"97e5cdc2",
   373 => x"32c84abf",
   374 => x"c27ea172",
   375 => x"6e48ebd9",
   376 => x"e6cdc278",
   377 => x"c848bf97",
   378 => x"d5c258a6",
   379 => x"c202bfde",
   380 => x"edc087cf",
   381 => x"c249bfe7",
   382 => x"714ae8ce",
   383 => x"e8e94bc8",
   384 => x"02987087",
   385 => x"c087c5c0",
   386 => x"87eac348",
   387 => x"bfd6d5c2",
   388 => x"ffd9c24c",
   389 => x"fbcdc25c",
   390 => x"c849bf97",
   391 => x"facdc231",
   392 => x"a14abf97",
   393 => x"fccdc249",
   394 => x"d04abf97",
   395 => x"49a17232",
   396 => x"97fdcdc2",
   397 => x"32d84abf",
   398 => x"c449a172",
   399 => x"d9c29166",
   400 => x"c281bfeb",
   401 => x"c259f3d9",
   402 => x"bf97c3ce",
   403 => x"c232c84a",
   404 => x"bf97c2ce",
   405 => x"c24aa24b",
   406 => x"bf97c4ce",
   407 => x"7333d04b",
   408 => x"cec24aa2",
   409 => x"4bbf97c5",
   410 => x"33d89bcf",
   411 => x"c24aa273",
   412 => x"c25af7d9",
   413 => x"c292748a",
   414 => x"7248f7d9",
   415 => x"c1c178a1",
   416 => x"e8cdc287",
   417 => x"c849bf97",
   418 => x"e7cdc231",
   419 => x"a14abf97",
   420 => x"c731c549",
   421 => x"29c981ff",
   422 => x"59ffd9c2",
   423 => x"97edcdc2",
   424 => x"32c84abf",
   425 => x"97eccdc2",
   426 => x"4aa24bbf",
   427 => x"6e9266c4",
   428 => x"fbd9c282",
   429 => x"f3d9c25a",
   430 => x"c278c048",
   431 => x"7248efd9",
   432 => x"d9c278a1",
   433 => x"d9c248ff",
   434 => x"c278bff3",
   435 => x"c248c3da",
   436 => x"78bff7d9",
   437 => x"bfded5c2",
   438 => x"87c9c002",
   439 => x"30c44874",
   440 => x"c9c07e70",
   441 => x"fbd9c287",
   442 => x"30c448bf",
   443 => x"d5c27e70",
   444 => x"786e48e2",
   445 => x"8ef848c1",
   446 => x"4c264d26",
   447 => x"4f264b26",
   448 => x"5c5b5e0e",
   449 => x"4a710e5d",
   450 => x"bfded5c2",
   451 => x"7287cb02",
   452 => x"722bc74b",
   453 => x"9dffc14d",
   454 => x"4b7287c9",
   455 => x"4d722bc8",
   456 => x"c29dffc3",
   457 => x"83bfebd9",
   458 => x"bfe3edc0",
   459 => x"87d902ab",
   460 => x"5be7edc0",
   461 => x"1ed6cdc2",
   462 => x"cbf14973",
   463 => x"7086c487",
   464 => x"87c50598",
   465 => x"e6c048c0",
   466 => x"ded5c287",
   467 => x"87d202bf",
   468 => x"91c44975",
   469 => x"81d6cdc2",
   470 => x"ffcf4c69",
   471 => x"9cffffff",
   472 => x"497587cb",
   473 => x"cdc291c2",
   474 => x"699f81d6",
   475 => x"fe48744c",
   476 => x"5e0e87c6",
   477 => x"0e5d5c5b",
   478 => x"4c7186f8",
   479 => x"87c5059c",
   480 => x"c1c348c0",
   481 => x"7ea4c887",
   482 => x"d878c048",
   483 => x"87c70266",
   484 => x"bf9766d8",
   485 => x"c087c505",
   486 => x"87eac248",
   487 => x"49c11ec0",
   488 => x"87e6c749",
   489 => x"4d7086c4",
   490 => x"c2c1029d",
   491 => x"e6d5c287",
   492 => x"4966d84a",
   493 => x"7087d7e2",
   494 => x"f2c00298",
   495 => x"d84a7587",
   496 => x"4bcb4966",
   497 => x"7087fce2",
   498 => x"e2c00298",
   499 => x"751ec087",
   500 => x"87c7029d",
   501 => x"c048a6c8",
   502 => x"c887c578",
   503 => x"78c148a6",
   504 => x"c64966c8",
   505 => x"86c487e4",
   506 => x"059d4d70",
   507 => x"7587fefe",
   508 => x"cfc1029d",
   509 => x"49a5dc87",
   510 => x"7869486e",
   511 => x"c449a5da",
   512 => x"a4c448a6",
   513 => x"48699f78",
   514 => x"780866c4",
   515 => x"bfded5c2",
   516 => x"d487d202",
   517 => x"699f49a5",
   518 => x"ffffc049",
   519 => x"d0487199",
   520 => x"c27e7030",
   521 => x"6e7ec087",
   522 => x"66c44849",
   523 => x"66c480bf",
   524 => x"7cc07808",
   525 => x"c449a4cc",
   526 => x"d079bf66",
   527 => x"79c049a4",
   528 => x"87c248c1",
   529 => x"8ef848c0",
   530 => x"0e87edfa",
   531 => x"5d5c5b5e",
   532 => x"9c4c710e",
   533 => x"87cbc102",
   534 => x"6949a4c8",
   535 => x"87c3c102",
   536 => x"6c4a66d0",
   537 => x"48a6d049",
   538 => x"4d78a172",
   539 => x"dad5c2b9",
   540 => x"baff4abf",
   541 => x"99719972",
   542 => x"87e4c002",
   543 => x"6b4ba4c4",
   544 => x"87fcf949",
   545 => x"d5c27b70",
   546 => x"6c49bfd6",
   547 => x"757c7181",
   548 => x"dad5c2b9",
   549 => x"baff4abf",
   550 => x"99719972",
   551 => x"87dcff05",
   552 => x"f97c66d0",
   553 => x"731e87d2",
   554 => x"9b4b711e",
   555 => x"c887c702",
   556 => x"056949a3",
   557 => x"48c087c5",
   558 => x"c287f6c0",
   559 => x"49bfefd9",
   560 => x"6a4aa3c4",
   561 => x"c28ac24a",
   562 => x"92bfd6d5",
   563 => x"c249a172",
   564 => x"4abfdad5",
   565 => x"a1729a6b",
   566 => x"e7edc049",
   567 => x"1e66c859",
   568 => x"87e4ea71",
   569 => x"987086c4",
   570 => x"c087c405",
   571 => x"c187c248",
   572 => x"87c8f848",
   573 => x"711e731e",
   574 => x"c0029b4b",
   575 => x"dac287e4",
   576 => x"4a735bc3",
   577 => x"d5c28ac2",
   578 => x"9249bfd6",
   579 => x"bfefd9c2",
   580 => x"c2807248",
   581 => x"7158c7da",
   582 => x"c230c448",
   583 => x"c058e6d5",
   584 => x"d9c287ed",
   585 => x"d9c248ff",
   586 => x"c278bff3",
   587 => x"c248c3da",
   588 => x"78bff7d9",
   589 => x"bfded5c2",
   590 => x"c287c902",
   591 => x"49bfd6d5",
   592 => x"87c731c4",
   593 => x"bffbd9c2",
   594 => x"c231c449",
   595 => x"f659e6d5",
   596 => x"5e0e87ea",
   597 => x"710e5c5b",
   598 => x"724bc04a",
   599 => x"e1c0029a",
   600 => x"49a2da87",
   601 => x"c24b699f",
   602 => x"02bfded5",
   603 => x"a2d487cf",
   604 => x"49699f49",
   605 => x"ffffc04c",
   606 => x"c234d09c",
   607 => x"744cc087",
   608 => x"4973b349",
   609 => x"f587edfd",
   610 => x"5e0e87f0",
   611 => x"0e5d5c5b",
   612 => x"4a7186f4",
   613 => x"9a727ec0",
   614 => x"c287d802",
   615 => x"c048d2cd",
   616 => x"cacdc278",
   617 => x"c3dac248",
   618 => x"cdc278bf",
   619 => x"d9c248ce",
   620 => x"c278bfff",
   621 => x"c048f3d5",
   622 => x"e2d5c250",
   623 => x"cdc249bf",
   624 => x"714abfd2",
   625 => x"c9c403aa",
   626 => x"cf497287",
   627 => x"e9c00599",
   628 => x"e3edc087",
   629 => x"cacdc248",
   630 => x"cdc278bf",
   631 => x"cdc21ed6",
   632 => x"c249bfca",
   633 => x"c148cacd",
   634 => x"e67178a1",
   635 => x"86c487da",
   636 => x"48dfedc0",
   637 => x"78d6cdc2",
   638 => x"edc087cc",
   639 => x"c048bfdf",
   640 => x"edc080e0",
   641 => x"cdc258e3",
   642 => x"c148bfd2",
   643 => x"d6cdc280",
   644 => x"0b5f2758",
   645 => x"97bf0000",
   646 => x"029d4dbf",
   647 => x"c387e3c2",
   648 => x"c202ade5",
   649 => x"edc087dc",
   650 => x"cb4bbfdf",
   651 => x"4c1149a3",
   652 => x"c105accf",
   653 => x"497587d2",
   654 => x"89c199df",
   655 => x"d5c291cd",
   656 => x"a3c181e6",
   657 => x"c351124a",
   658 => x"51124aa3",
   659 => x"124aa3c5",
   660 => x"4aa3c751",
   661 => x"a3c95112",
   662 => x"ce51124a",
   663 => x"51124aa3",
   664 => x"124aa3d0",
   665 => x"4aa3d251",
   666 => x"a3d45112",
   667 => x"d651124a",
   668 => x"51124aa3",
   669 => x"124aa3d8",
   670 => x"4aa3dc51",
   671 => x"a3de5112",
   672 => x"c151124a",
   673 => x"87fac07e",
   674 => x"99c84974",
   675 => x"87ebc005",
   676 => x"99d04974",
   677 => x"dc87d105",
   678 => x"cbc00266",
   679 => x"dc497387",
   680 => x"98700f66",
   681 => x"87d3c002",
   682 => x"c6c0056e",
   683 => x"e6d5c287",
   684 => x"c050c048",
   685 => x"48bfdfed",
   686 => x"c287dfc2",
   687 => x"c048f3d5",
   688 => x"d5c27e50",
   689 => x"c249bfe2",
   690 => x"4abfd2cd",
   691 => x"fb04aa71",
   692 => x"dac287f7",
   693 => x"c005bfc3",
   694 => x"d5c287c8",
   695 => x"c102bfde",
   696 => x"cdc287f6",
   697 => x"f049bfce",
   698 => x"cdc287d6",
   699 => x"a6c458d2",
   700 => x"cecdc248",
   701 => x"d5c278bf",
   702 => x"c002bfde",
   703 => x"66c487d8",
   704 => x"ffffcf49",
   705 => x"a999f8ff",
   706 => x"87c5c002",
   707 => x"e1c04cc0",
   708 => x"c04cc187",
   709 => x"66c487dc",
   710 => x"f8ffcf49",
   711 => x"c002a999",
   712 => x"a6c887c8",
   713 => x"c078c048",
   714 => x"a6c887c5",
   715 => x"c878c148",
   716 => x"9c744c66",
   717 => x"87e0c005",
   718 => x"c24966c4",
   719 => x"d6d5c289",
   720 => x"c2914abf",
   721 => x"4abfefd9",
   722 => x"48cacdc2",
   723 => x"c278a172",
   724 => x"c048d2cd",
   725 => x"87e1f978",
   726 => x"8ef448c0",
   727 => x"0087d9ee",
   728 => x"ff000000",
   729 => x"6fffffff",
   730 => x"7800000b",
   731 => x"4600000b",
   732 => x"32335441",
   733 => x"00202020",
   734 => x"31544146",
   735 => x"20202036",
   736 => x"d4ff1e00",
   737 => x"78ffc348",
   738 => x"4f264868",
   739 => x"48d4ff1e",
   740 => x"ff78ffc3",
   741 => x"e1c048d0",
   742 => x"48d4ff78",
   743 => x"dac278d4",
   744 => x"d4ff48c7",
   745 => x"4f2650bf",
   746 => x"48d0ff1e",
   747 => x"2678e0c0",
   748 => x"ccff1e4f",
   749 => x"99497087",
   750 => x"c087c602",
   751 => x"f105a9fb",
   752 => x"26487187",
   753 => x"5b5e0e4f",
   754 => x"4b710e5c",
   755 => x"f0fe4cc0",
   756 => x"99497087",
   757 => x"87f9c002",
   758 => x"02a9ecc0",
   759 => x"c087f2c0",
   760 => x"c002a9fb",
   761 => x"66cc87eb",
   762 => x"c703acb7",
   763 => x"0266d087",
   764 => x"537187c2",
   765 => x"c2029971",
   766 => x"fe84c187",
   767 => x"497087c3",
   768 => x"87cd0299",
   769 => x"02a9ecc0",
   770 => x"fbc087c7",
   771 => x"d5ff05a9",
   772 => x"0266d087",
   773 => x"97c087c3",
   774 => x"a9ecc07b",
   775 => x"7487c405",
   776 => x"7487c54a",
   777 => x"8a0ac04a",
   778 => x"87c24872",
   779 => x"4c264d26",
   780 => x"4f264b26",
   781 => x"87c9fd1e",
   782 => x"f0c04a70",
   783 => x"87c904aa",
   784 => x"01aaf9c0",
   785 => x"f0c087c3",
   786 => x"aac1c18a",
   787 => x"c187c904",
   788 => x"c301aada",
   789 => x"8af7c087",
   790 => x"4f264872",
   791 => x"5c5b5e0e",
   792 => x"86f80e5d",
   793 => x"4dc04c71",
   794 => x"c087e1fc",
   795 => x"fbf3c04b",
   796 => x"c049bf97",
   797 => x"87cf04a9",
   798 => x"c187f6fc",
   799 => x"fbf3c083",
   800 => x"ab49bf97",
   801 => x"c087f106",
   802 => x"bf97fbf3",
   803 => x"fb87cf02",
   804 => x"497087ef",
   805 => x"87c60299",
   806 => x"05a9ecc0",
   807 => x"4bc087f1",
   808 => x"7087defb",
   809 => x"87d9fb7e",
   810 => x"fb58a6c8",
   811 => x"4a7087d3",
   812 => x"a4c883c1",
   813 => x"49699749",
   814 => x"da05a96e",
   815 => x"49a4c987",
   816 => x"c4496997",
   817 => x"ce05a966",
   818 => x"49a4ca87",
   819 => x"aa496997",
   820 => x"c187c405",
   821 => x"6e87d44d",
   822 => x"a8ecc048",
   823 => x"6e87c802",
   824 => x"a8fbc048",
   825 => x"c087c405",
   826 => x"754dc14b",
   827 => x"effe029d",
   828 => x"87f4fa87",
   829 => x"8ef84873",
   830 => x"0087f1fc",
   831 => x"5c5b5e0e",
   832 => x"86f80e5d",
   833 => x"d4ff7e71",
   834 => x"c21e6e4b",
   835 => x"e949ccda",
   836 => x"86c487e0",
   837 => x"c4029870",
   838 => x"ddc187ea",
   839 => x"6e4dbfe2",
   840 => x"87f8fc49",
   841 => x"7058a6c8",
   842 => x"87c50598",
   843 => x"c148a6c4",
   844 => x"48d0ff78",
   845 => x"d5c178c5",
   846 => x"4966c47b",
   847 => x"31c689c1",
   848 => x"97e0ddc1",
   849 => x"71484abf",
   850 => x"ff7b70b0",
   851 => x"78c448d0",
   852 => x"97c7dac2",
   853 => x"99d049bf",
   854 => x"c587d702",
   855 => x"7bd6c178",
   856 => x"ffc34ac0",
   857 => x"c082c17b",
   858 => x"f504aae0",
   859 => x"48d0ff87",
   860 => x"ffc378c4",
   861 => x"48d0ff7b",
   862 => x"d3c178c5",
   863 => x"c47bc17b",
   864 => x"adb7c078",
   865 => x"87ebc206",
   866 => x"bfd4dac2",
   867 => x"029c8d4c",
   868 => x"c287c2c2",
   869 => x"c47ed6cd",
   870 => x"c0c848a6",
   871 => x"b7c08c78",
   872 => x"87c603ac",
   873 => x"78a4c0c8",
   874 => x"dac24cc0",
   875 => x"49bf97c7",
   876 => x"d00299d0",
   877 => x"c21ec087",
   878 => x"eb49ccda",
   879 => x"86c487e8",
   880 => x"f5c04a70",
   881 => x"d6cdc287",
   882 => x"ccdac21e",
   883 => x"87d6eb49",
   884 => x"4a7086c4",
   885 => x"c848d0ff",
   886 => x"d4c178c5",
   887 => x"bf976e7b",
   888 => x"c1486e7b",
   889 => x"c47e7080",
   890 => x"88c14866",
   891 => x"7058a6c8",
   892 => x"e8ff0598",
   893 => x"48d0ff87",
   894 => x"9a7278c4",
   895 => x"c087c505",
   896 => x"87c2c148",
   897 => x"dac21ec1",
   898 => x"fee849cc",
   899 => x"7486c487",
   900 => x"fefd059c",
   901 => x"adb7c087",
   902 => x"c287d106",
   903 => x"c048ccda",
   904 => x"c080d078",
   905 => x"c280f478",
   906 => x"78bfd8da",
   907 => x"01adb7c0",
   908 => x"ff87d5fd",
   909 => x"78c548d0",
   910 => x"c07bd3c1",
   911 => x"c178c47b",
   912 => x"87c2c048",
   913 => x"8ef848c0",
   914 => x"4c264d26",
   915 => x"4f264b26",
   916 => x"5c5b5e0e",
   917 => x"711e0e5d",
   918 => x"4d4cc04b",
   919 => x"e8c004ab",
   920 => x"dcf1c087",
   921 => x"029d751e",
   922 => x"4ac087c4",
   923 => x"4ac187c2",
   924 => x"d5ec4972",
   925 => x"7086c487",
   926 => x"6e84c17e",
   927 => x"7387c205",
   928 => x"7385c14c",
   929 => x"d8ff06ac",
   930 => x"26486e87",
   931 => x"1e87f9fe",
   932 => x"66c44a71",
   933 => x"7287c505",
   934 => x"87e0f949",
   935 => x"5e0e4f26",
   936 => x"0e5d5c5b",
   937 => x"494c711e",
   938 => x"dac291de",
   939 => x"85714df4",
   940 => x"c1026d97",
   941 => x"dac287dc",
   942 => x"7449bfe0",
   943 => x"cffe7181",
   944 => x"487e7087",
   945 => x"f2c00298",
   946 => x"e8dac287",
   947 => x"cb4a704b",
   948 => x"d2c7ff49",
   949 => x"cb4b7487",
   950 => x"f4ddc193",
   951 => x"c083c483",
   952 => x"747bd6fc",
   953 => x"ecc0c149",
   954 => x"c17b7587",
   955 => x"bf97e1dd",
   956 => x"dac21e49",
   957 => x"d6fe49e8",
   958 => x"7486c487",
   959 => x"d4c0c149",
   960 => x"c149c087",
   961 => x"c287f3c1",
   962 => x"c048c8da",
   963 => x"dd49c178",
   964 => x"fc2687f9",
   965 => x"6f4c87f2",
   966 => x"6e696461",
   967 => x"2e2e2e67",
   968 => x"1e731e00",
   969 => x"c2494a71",
   970 => x"81bfe0da",
   971 => x"87e0fc71",
   972 => x"029b4b70",
   973 => x"e84987c4",
   974 => x"dac287d8",
   975 => x"78c048e0",
   976 => x"c6dd49c1",
   977 => x"87c4fc87",
   978 => x"c149c01e",
   979 => x"2687ebc0",
   980 => x"4a711e4f",
   981 => x"c191cb49",
   982 => x"c881f4dd",
   983 => x"c2481181",
   984 => x"c258ccda",
   985 => x"c048e0da",
   986 => x"dc49c178",
   987 => x"4f2687dd",
   988 => x"0299711e",
   989 => x"dfc187d2",
   990 => x"50c048c9",
   991 => x"fdc080f7",
   992 => x"ddc140d1",
   993 => x"87ce78ed",
   994 => x"48c5dfc1",
   995 => x"78e6ddc1",
   996 => x"fdc080fc",
   997 => x"4f2678c8",
   998 => x"5c5b5e0e",
   999 => x"86f40e5d",
  1000 => x"4dd6cdc2",
  1001 => x"a6c44cc0",
  1002 => x"c278c048",
  1003 => x"48bfe0da",
  1004 => x"c106a8c0",
  1005 => x"cdc287c0",
  1006 => x"029848d6",
  1007 => x"c087f7c0",
  1008 => x"c81edcf1",
  1009 => x"87c70266",
  1010 => x"c048a6c4",
  1011 => x"c487c578",
  1012 => x"78c148a6",
  1013 => x"e64966c4",
  1014 => x"86c487f0",
  1015 => x"84c14d70",
  1016 => x"c14866c4",
  1017 => x"58a6c880",
  1018 => x"bfe0dac2",
  1019 => x"87c603ac",
  1020 => x"ff059d75",
  1021 => x"4cc087c9",
  1022 => x"c3029d75",
  1023 => x"f1c087dc",
  1024 => x"66c81edc",
  1025 => x"cc87c702",
  1026 => x"78c048a6",
  1027 => x"a6cc87c5",
  1028 => x"cc78c148",
  1029 => x"f1e54966",
  1030 => x"7086c487",
  1031 => x"0298487e",
  1032 => x"4987e4c2",
  1033 => x"699781cb",
  1034 => x"0299d049",
  1035 => x"7487d4c1",
  1036 => x"c191cb49",
  1037 => x"c081f4dd",
  1038 => x"c879e1fc",
  1039 => x"51ffc381",
  1040 => x"91de4974",
  1041 => x"4df4dac2",
  1042 => x"c1c28571",
  1043 => x"a5c17d97",
  1044 => x"51e0c049",
  1045 => x"97e6d5c2",
  1046 => x"87d202bf",
  1047 => x"a5c284c1",
  1048 => x"e6d5c24b",
  1049 => x"ff49db4a",
  1050 => x"c187fcc0",
  1051 => x"a5cd87d9",
  1052 => x"c151c049",
  1053 => x"4ba5c284",
  1054 => x"49cb4a6e",
  1055 => x"87e7c0ff",
  1056 => x"7487c4c1",
  1057 => x"c191cb49",
  1058 => x"c081f4dd",
  1059 => x"c279defa",
  1060 => x"bf97e6d5",
  1061 => x"7487d802",
  1062 => x"c191de49",
  1063 => x"f4dac284",
  1064 => x"c283714b",
  1065 => x"dd4ae6d5",
  1066 => x"fafffe49",
  1067 => x"7487d887",
  1068 => x"c293de4b",
  1069 => x"cb83f4da",
  1070 => x"51c049a3",
  1071 => x"6e7384c1",
  1072 => x"fe49cb4a",
  1073 => x"c487e0ff",
  1074 => x"80c14866",
  1075 => x"c758a6c8",
  1076 => x"c5c003ac",
  1077 => x"fc056e87",
  1078 => x"487487e4",
  1079 => x"e7f58ef4",
  1080 => x"1e731e87",
  1081 => x"cb494b71",
  1082 => x"f4ddc191",
  1083 => x"4aa1c881",
  1084 => x"48e0ddc1",
  1085 => x"a1c95012",
  1086 => x"fbf3c04a",
  1087 => x"ca501248",
  1088 => x"e1ddc181",
  1089 => x"c1501148",
  1090 => x"bf97e1dd",
  1091 => x"49c01e49",
  1092 => x"c287fcf5",
  1093 => x"de48c8da",
  1094 => x"d549c178",
  1095 => x"f42687ed",
  1096 => x"5e0e87ea",
  1097 => x"0e5d5c5b",
  1098 => x"4d7186f4",
  1099 => x"c191cb49",
  1100 => x"c881f4dd",
  1101 => x"a1ca4aa1",
  1102 => x"48a6c47e",
  1103 => x"bfd0dec2",
  1104 => x"bf976e78",
  1105 => x"4c66c44b",
  1106 => x"48122c73",
  1107 => x"7058a6cc",
  1108 => x"c984c19c",
  1109 => x"49699781",
  1110 => x"c204acb7",
  1111 => x"6e4cc087",
  1112 => x"c84abf97",
  1113 => x"31724966",
  1114 => x"66c4b9ff",
  1115 => x"72487499",
  1116 => x"484a7030",
  1117 => x"dec2b071",
  1118 => x"e4c058d4",
  1119 => x"49c087d7",
  1120 => x"7587c8d4",
  1121 => x"ccf6c049",
  1122 => x"f28ef487",
  1123 => x"731e87fa",
  1124 => x"494b711e",
  1125 => x"7387cbfe",
  1126 => x"87c6fe49",
  1127 => x"1e87edf2",
  1128 => x"4b711e73",
  1129 => x"024aa3c6",
  1130 => x"8ac187db",
  1131 => x"8a87d602",
  1132 => x"87dac102",
  1133 => x"fcc0028a",
  1134 => x"c0028a87",
  1135 => x"028a87e1",
  1136 => x"dbc187cb",
  1137 => x"f649c787",
  1138 => x"dec187c7",
  1139 => x"e0dac287",
  1140 => x"cbc102bf",
  1141 => x"88c14887",
  1142 => x"58e4dac2",
  1143 => x"c287c1c1",
  1144 => x"02bfe4da",
  1145 => x"c287f9c0",
  1146 => x"48bfe0da",
  1147 => x"dac280c1",
  1148 => x"ebc058e4",
  1149 => x"e0dac287",
  1150 => x"89c649bf",
  1151 => x"59e4dac2",
  1152 => x"03a9b7c0",
  1153 => x"dac287da",
  1154 => x"78c048e0",
  1155 => x"dac287d2",
  1156 => x"cb02bfe4",
  1157 => x"e0dac287",
  1158 => x"80c648bf",
  1159 => x"58e4dac2",
  1160 => x"e6d149c0",
  1161 => x"c0497387",
  1162 => x"f087eaf3",
  1163 => x"5e0e87de",
  1164 => x"0e5d5c5b",
  1165 => x"dc86d4ff",
  1166 => x"a6c859a6",
  1167 => x"c478c048",
  1168 => x"66c0c180",
  1169 => x"c180c478",
  1170 => x"c180c478",
  1171 => x"e4dac278",
  1172 => x"c278c148",
  1173 => x"48bfc8da",
  1174 => x"c905a8de",
  1175 => x"87f8f487",
  1176 => x"cf58a6cc",
  1177 => x"e3e487e4",
  1178 => x"87c5e587",
  1179 => x"7087d2e4",
  1180 => x"acfbc04c",
  1181 => x"87fbc102",
  1182 => x"c10566d8",
  1183 => x"fcc087ed",
  1184 => x"82c44a66",
  1185 => x"1e727e6a",
  1186 => x"48ffd9c1",
  1187 => x"c84966c4",
  1188 => x"41204aa1",
  1189 => x"f905aa71",
  1190 => x"26511087",
  1191 => x"66fcc04a",
  1192 => x"e1c3c148",
  1193 => x"c7496a78",
  1194 => x"c0517481",
  1195 => x"c84966fc",
  1196 => x"c051c181",
  1197 => x"c94966fc",
  1198 => x"c051c081",
  1199 => x"ca4966fc",
  1200 => x"c151c081",
  1201 => x"6a1ed81e",
  1202 => x"e381c849",
  1203 => x"86c887f7",
  1204 => x"4866c0c1",
  1205 => x"c701a8c0",
  1206 => x"48a6c887",
  1207 => x"87ce78c1",
  1208 => x"4866c0c1",
  1209 => x"a6d088c1",
  1210 => x"e387c358",
  1211 => x"a6d087c3",
  1212 => x"7478c248",
  1213 => x"cdcd029c",
  1214 => x"4866c887",
  1215 => x"a866c4c1",
  1216 => x"87c2cd03",
  1217 => x"c048a6dc",
  1218 => x"c080e878",
  1219 => x"87f1e178",
  1220 => x"d0c14c70",
  1221 => x"d5c205ac",
  1222 => x"7e66c487",
  1223 => x"c887d5e4",
  1224 => x"dce158a6",
  1225 => x"c04c7087",
  1226 => x"c105acec",
  1227 => x"66c887eb",
  1228 => x"c091cb49",
  1229 => x"c48166fc",
  1230 => x"4d6a4aa1",
  1231 => x"c44aa1c8",
  1232 => x"fdc05266",
  1233 => x"f8e079d1",
  1234 => x"9c4c7087",
  1235 => x"c087d802",
  1236 => x"d202acfb",
  1237 => x"e0557487",
  1238 => x"4c7087e7",
  1239 => x"87c7029c",
  1240 => x"05acfbc0",
  1241 => x"c087eeff",
  1242 => x"c1c255e0",
  1243 => x"7d97c055",
  1244 => x"6e4866d8",
  1245 => x"87db05a8",
  1246 => x"cc4866c8",
  1247 => x"ca04a866",
  1248 => x"4866c887",
  1249 => x"a6cc80c1",
  1250 => x"cc87c858",
  1251 => x"88c14866",
  1252 => x"ff58a6d0",
  1253 => x"7087eadf",
  1254 => x"acd0c14c",
  1255 => x"d487c805",
  1256 => x"80c14866",
  1257 => x"c158a6d8",
  1258 => x"fd02acd0",
  1259 => x"66c487eb",
  1260 => x"a866d848",
  1261 => x"87e0c905",
  1262 => x"48a6e0c0",
  1263 => x"487478c0",
  1264 => x"7088fbc0",
  1265 => x"0298487e",
  1266 => x"4887e2c9",
  1267 => x"7e7088cb",
  1268 => x"c1029848",
  1269 => x"c94887cd",
  1270 => x"487e7088",
  1271 => x"fec30298",
  1272 => x"88c44887",
  1273 => x"98487e70",
  1274 => x"4887ce02",
  1275 => x"7e7088c1",
  1276 => x"c3029848",
  1277 => x"d6c887e9",
  1278 => x"48a6dc87",
  1279 => x"ff78f0c0",
  1280 => x"7087fedd",
  1281 => x"acecc04c",
  1282 => x"87c4c002",
  1283 => x"5ca6e0c0",
  1284 => x"02acecc0",
  1285 => x"ddff87cd",
  1286 => x"4c7087e7",
  1287 => x"05acecc0",
  1288 => x"c087f3ff",
  1289 => x"c002acec",
  1290 => x"ddff87c4",
  1291 => x"1ec087d3",
  1292 => x"66d01eca",
  1293 => x"c191cb49",
  1294 => x"714866c4",
  1295 => x"58a6cc80",
  1296 => x"c44866c8",
  1297 => x"58a6d080",
  1298 => x"49bf66cc",
  1299 => x"87f5ddff",
  1300 => x"1ede1ec1",
  1301 => x"49bf66d4",
  1302 => x"87e9ddff",
  1303 => x"497086d0",
  1304 => x"8808c048",
  1305 => x"58a6e8c0",
  1306 => x"c006a8c0",
  1307 => x"e4c087ee",
  1308 => x"a8dd4866",
  1309 => x"87e4c003",
  1310 => x"49bf66c4",
  1311 => x"8166e4c0",
  1312 => x"c051e0c0",
  1313 => x"c14966e4",
  1314 => x"bf66c481",
  1315 => x"51c1c281",
  1316 => x"4966e4c0",
  1317 => x"66c481c2",
  1318 => x"51c081bf",
  1319 => x"c3c1486e",
  1320 => x"496e78e1",
  1321 => x"66d081c8",
  1322 => x"c9496e51",
  1323 => x"5166d481",
  1324 => x"81ca496e",
  1325 => x"d05166dc",
  1326 => x"80c14866",
  1327 => x"c858a6d4",
  1328 => x"66cc4866",
  1329 => x"cbc004a8",
  1330 => x"4866c887",
  1331 => x"a6cc80c1",
  1332 => x"87d9c558",
  1333 => x"c14866cc",
  1334 => x"58a6d088",
  1335 => x"ff87cec5",
  1336 => x"c087d1dd",
  1337 => x"ff58a6e8",
  1338 => x"c087c9dd",
  1339 => x"c058a6e0",
  1340 => x"c005a8ec",
  1341 => x"a6dc87ca",
  1342 => x"66e4c048",
  1343 => x"87c4c078",
  1344 => x"87fdd9ff",
  1345 => x"cb4966c8",
  1346 => x"66fcc091",
  1347 => x"70807148",
  1348 => x"82c84a7e",
  1349 => x"81ca496e",
  1350 => x"5166e4c0",
  1351 => x"c14966dc",
  1352 => x"66e4c081",
  1353 => x"7148c189",
  1354 => x"c1497030",
  1355 => x"7a977189",
  1356 => x"bfd0dec2",
  1357 => x"66e4c049",
  1358 => x"4a6a9729",
  1359 => x"c0987148",
  1360 => x"6e58a6ec",
  1361 => x"6981c449",
  1362 => x"4866d84d",
  1363 => x"02a866c4",
  1364 => x"c487c8c0",
  1365 => x"78c048a6",
  1366 => x"c487c5c0",
  1367 => x"78c148a6",
  1368 => x"c01e66c4",
  1369 => x"49751ee0",
  1370 => x"87d9d9ff",
  1371 => x"4c7086c8",
  1372 => x"06acb7c0",
  1373 => x"7487d4c1",
  1374 => x"49e0c085",
  1375 => x"4b758974",
  1376 => x"4ac8dac1",
  1377 => x"deecfe71",
  1378 => x"c085c287",
  1379 => x"c14866e0",
  1380 => x"a6e4c080",
  1381 => x"66e8c058",
  1382 => x"7081c149",
  1383 => x"c8c002a9",
  1384 => x"48a6c487",
  1385 => x"c5c078c0",
  1386 => x"48a6c487",
  1387 => x"66c478c1",
  1388 => x"49a4c21e",
  1389 => x"7148e0c0",
  1390 => x"1e497088",
  1391 => x"d8ff4975",
  1392 => x"86c887c3",
  1393 => x"01a8b7c0",
  1394 => x"c087c0ff",
  1395 => x"c00266e0",
  1396 => x"496e87d1",
  1397 => x"e0c081c9",
  1398 => x"486e5166",
  1399 => x"78e2c4c1",
  1400 => x"6e87ccc0",
  1401 => x"c281c949",
  1402 => x"c1486e51",
  1403 => x"c878cec6",
  1404 => x"66cc4866",
  1405 => x"cbc004a8",
  1406 => x"4866c887",
  1407 => x"a6cc80c1",
  1408 => x"87e9c058",
  1409 => x"c14866cc",
  1410 => x"58a6d088",
  1411 => x"ff87dec0",
  1412 => x"7087ded6",
  1413 => x"87d5c04c",
  1414 => x"05acc6c1",
  1415 => x"d087c8c0",
  1416 => x"80c14866",
  1417 => x"ff58a6d4",
  1418 => x"7087c6d6",
  1419 => x"4866d44c",
  1420 => x"a6d880c1",
  1421 => x"029c7458",
  1422 => x"c887cbc0",
  1423 => x"c4c14866",
  1424 => x"f204a866",
  1425 => x"d5ff87fe",
  1426 => x"66c887de",
  1427 => x"03a8c748",
  1428 => x"c287e5c0",
  1429 => x"c048e4da",
  1430 => x"4966c878",
  1431 => x"fcc091cb",
  1432 => x"a1c48166",
  1433 => x"c04a6a4a",
  1434 => x"66c87952",
  1435 => x"cc80c148",
  1436 => x"a8c758a6",
  1437 => x"87dbff04",
  1438 => x"ff8ed4ff",
  1439 => x"4c87c9df",
  1440 => x"2064616f",
  1441 => x"00202e2a",
  1442 => x"1e00203a",
  1443 => x"4b711e73",
  1444 => x"87c6029b",
  1445 => x"48e0dac2",
  1446 => x"1ec778c0",
  1447 => x"bfe0dac2",
  1448 => x"f4ddc11e",
  1449 => x"c8dac21e",
  1450 => x"c1ee49bf",
  1451 => x"c286cc87",
  1452 => x"49bfc8da",
  1453 => x"7387f9e2",
  1454 => x"87c8029b",
  1455 => x"49f4ddc1",
  1456 => x"87e3e2c0",
  1457 => x"87c4deff",
  1458 => x"e0ddc11e",
  1459 => x"c150c048",
  1460 => x"49bfd7df",
  1461 => x"87e4d8ff",
  1462 => x"4f2648c0",
  1463 => x"87dec71e",
  1464 => x"e6fe49c1",
  1465 => x"c7effe87",
  1466 => x"02987087",
  1467 => x"f6fe87cd",
  1468 => x"987087e1",
  1469 => x"c187c402",
  1470 => x"c087c24a",
  1471 => x"059a724a",
  1472 => x"1ec087ce",
  1473 => x"49f7dcc1",
  1474 => x"87deeec0",
  1475 => x"87fe86c4",
  1476 => x"48e0dac2",
  1477 => x"dac278c0",
  1478 => x"78c048c8",
  1479 => x"c2ddc11e",
  1480 => x"c5eec049",
  1481 => x"fe1ec087",
  1482 => x"497087de",
  1483 => x"87faedc0",
  1484 => x"f887cac3",
  1485 => x"534f268e",
  1486 => x"61662044",
  1487 => x"64656c69",
  1488 => x"6f42002e",
  1489 => x"6e69746f",
  1490 => x"2e2e2e67",
  1491 => x"e2c01e00",
  1492 => x"87fa87d2",
  1493 => x"fe1e4f26",
  1494 => x"87f187c2",
  1495 => x"4f2648c0",
  1496 => x"00010000",
  1497 => x"20800000",
  1498 => x"74697845",
  1499 => x"42208000",
  1500 => x"006b6361",
  1501 => x"00000e9e",
  1502 => x"000026b4",
  1503 => x"9e000000",
  1504 => x"d200000e",
  1505 => x"00000026",
  1506 => x"0e9e0000",
  1507 => x"26f00000",
  1508 => x"00000000",
  1509 => x"000e9e00",
  1510 => x"00270e00",
  1511 => x"00000000",
  1512 => x"00000e9e",
  1513 => x"0000272c",
  1514 => x"9e000000",
  1515 => x"4a00000e",
  1516 => x"00000027",
  1517 => x"0e9e0000",
  1518 => x"27680000",
  1519 => x"00000000",
  1520 => x"000f5100",
  1521 => x"00000000",
  1522 => x"00000000",
  1523 => x"0000119f",
  1524 => x"00000000",
  1525 => x"db000000",
  1526 => x"42000017",
  1527 => x"20544f4f",
  1528 => x"52202020",
  1529 => x"1e004d4f",
  1530 => x"c048f0fe",
  1531 => x"7909cd78",
  1532 => x"1e4f2609",
  1533 => x"bff0fe1e",
  1534 => x"2626487e",
  1535 => x"f0fe1e4f",
  1536 => x"2678c148",
  1537 => x"f0fe1e4f",
  1538 => x"2678c048",
  1539 => x"4a711e4f",
  1540 => x"265252c0",
  1541 => x"5b5e0e4f",
  1542 => x"f40e5d5c",
  1543 => x"974d7186",
  1544 => x"a5c17e6d",
  1545 => x"486c974c",
  1546 => x"6e58a6c8",
  1547 => x"a866c448",
  1548 => x"ff87c505",
  1549 => x"87e6c048",
  1550 => x"c287caff",
  1551 => x"6c9749a5",
  1552 => x"4ba3714b",
  1553 => x"974b6b97",
  1554 => x"486e7e6c",
  1555 => x"a6c880c1",
  1556 => x"cc98c758",
  1557 => x"977058a6",
  1558 => x"87e1fe7c",
  1559 => x"8ef44873",
  1560 => x"4c264d26",
  1561 => x"4f264b26",
  1562 => x"5c5b5e0e",
  1563 => x"7186f40e",
  1564 => x"4a66d84c",
  1565 => x"c29affc3",
  1566 => x"6c974ba4",
  1567 => x"49a17349",
  1568 => x"6c975172",
  1569 => x"c1486e7e",
  1570 => x"58a6c880",
  1571 => x"a6cc98c7",
  1572 => x"f4547058",
  1573 => x"87caff8e",
  1574 => x"e8fd1e1e",
  1575 => x"4abfe087",
  1576 => x"c0e0c049",
  1577 => x"87cb0299",
  1578 => x"dec21e72",
  1579 => x"f7fe49c6",
  1580 => x"fc86c487",
  1581 => x"7e7087fd",
  1582 => x"2687c2fd",
  1583 => x"c21e4f26",
  1584 => x"fd49c6de",
  1585 => x"e2c187c7",
  1586 => x"dafc49d8",
  1587 => x"87eec387",
  1588 => x"5e0e4f26",
  1589 => x"0e5d5c5b",
  1590 => x"dec24d71",
  1591 => x"f4fc49c6",
  1592 => x"c04b7087",
  1593 => x"c304abb7",
  1594 => x"f0c387c2",
  1595 => x"87c905ab",
  1596 => x"48f6e6c1",
  1597 => x"e3c278c1",
  1598 => x"abe0c387",
  1599 => x"c187c905",
  1600 => x"c148fae6",
  1601 => x"87d4c278",
  1602 => x"bffae6c1",
  1603 => x"c287c602",
  1604 => x"c24ca3c0",
  1605 => x"c14c7387",
  1606 => x"02bff6e6",
  1607 => x"7487e0c0",
  1608 => x"29b7c449",
  1609 => x"cde8c191",
  1610 => x"cf4a7481",
  1611 => x"c192c29a",
  1612 => x"70307248",
  1613 => x"72baff4a",
  1614 => x"70986948",
  1615 => x"7487db79",
  1616 => x"29b7c449",
  1617 => x"cde8c191",
  1618 => x"cf4a7481",
  1619 => x"c392c29a",
  1620 => x"70307248",
  1621 => x"b069484a",
  1622 => x"9d757970",
  1623 => x"87f0c005",
  1624 => x"c848d0ff",
  1625 => x"d4ff78e1",
  1626 => x"c178c548",
  1627 => x"02bffae6",
  1628 => x"e0c387c3",
  1629 => x"f6e6c178",
  1630 => x"87c602bf",
  1631 => x"c348d4ff",
  1632 => x"d4ff78f0",
  1633 => x"ff0b7b0b",
  1634 => x"e1c848d0",
  1635 => x"78e0c078",
  1636 => x"48fae6c1",
  1637 => x"e6c178c0",
  1638 => x"78c048f6",
  1639 => x"49c6dec2",
  1640 => x"7087f2f9",
  1641 => x"abb7c04b",
  1642 => x"87fefc03",
  1643 => x"4d2648c0",
  1644 => x"4b264c26",
  1645 => x"00004f26",
  1646 => x"00000000",
  1647 => x"c01e0000",
  1648 => x"c449724a",
  1649 => x"cde8c191",
  1650 => x"c179c081",
  1651 => x"aab7d082",
  1652 => x"2687ee04",
  1653 => x"5b5e0e4f",
  1654 => x"710e5d5c",
  1655 => x"87e5f84d",
  1656 => x"b7c44a75",
  1657 => x"e8c1922a",
  1658 => x"4c7582cd",
  1659 => x"94c29ccf",
  1660 => x"744b496a",
  1661 => x"c29bc32b",
  1662 => x"70307448",
  1663 => x"74bcff4c",
  1664 => x"70987148",
  1665 => x"87f5f77a",
  1666 => x"e1fe4873",
  1667 => x"00000087",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"d0ff1e00",
  1684 => x"78e1c848",
  1685 => x"d4ff4871",
  1686 => x"66c47808",
  1687 => x"08d4ff48",
  1688 => x"1e4f2678",
  1689 => x"66c44a71",
  1690 => x"49721e49",
  1691 => x"ff87deff",
  1692 => x"e0c048d0",
  1693 => x"4f262678",
  1694 => x"711e731e",
  1695 => x"4966c84b",
  1696 => x"c14a731e",
  1697 => x"ff49a2e0",
  1698 => x"c42687d9",
  1699 => x"264d2687",
  1700 => x"264b264c",
  1701 => x"d4ff1e4f",
  1702 => x"7affc34a",
  1703 => x"c048d0ff",
  1704 => x"7ade78e1",
  1705 => x"bfd0dec2",
  1706 => x"c848497a",
  1707 => x"717a7028",
  1708 => x"7028d048",
  1709 => x"d848717a",
  1710 => x"ff7a7028",
  1711 => x"e0c048d0",
  1712 => x"1e4f2678",
  1713 => x"c848d0ff",
  1714 => x"487178c9",
  1715 => x"7808d4ff",
  1716 => x"711e4f26",
  1717 => x"87eb494a",
  1718 => x"c848d0ff",
  1719 => x"1e4f2678",
  1720 => x"4b711e73",
  1721 => x"bfe0dec2",
  1722 => x"c287c302",
  1723 => x"d0ff87eb",
  1724 => x"78c9c848",
  1725 => x"e0c04873",
  1726 => x"08d4ffb0",
  1727 => x"d4dec278",
  1728 => x"c878c048",
  1729 => x"87c50266",
  1730 => x"c249ffc3",
  1731 => x"c249c087",
  1732 => x"cc59dcde",
  1733 => x"87c60266",
  1734 => x"4ad5d5c5",
  1735 => x"ffcf87c4",
  1736 => x"dec24aff",
  1737 => x"dec25ae0",
  1738 => x"78c148e0",
  1739 => x"4d2687c4",
  1740 => x"4b264c26",
  1741 => x"5e0e4f26",
  1742 => x"0e5d5c5b",
  1743 => x"dec24a71",
  1744 => x"724cbfdc",
  1745 => x"87cb029a",
  1746 => x"c191c849",
  1747 => x"714bd5eb",
  1748 => x"c187c483",
  1749 => x"c04bd5ef",
  1750 => x"7449134d",
  1751 => x"d8dec299",
  1752 => x"b87148bf",
  1753 => x"7808d4ff",
  1754 => x"852cb7c1",
  1755 => x"04adb7c8",
  1756 => x"dec287e7",
  1757 => x"c848bfd4",
  1758 => x"d8dec280",
  1759 => x"87eefe58",
  1760 => x"711e731e",
  1761 => x"9a4a134b",
  1762 => x"7287cb02",
  1763 => x"87e6fe49",
  1764 => x"059a4a13",
  1765 => x"d9fe87f5",
  1766 => x"dec21e87",
  1767 => x"c249bfd4",
  1768 => x"c148d4de",
  1769 => x"c0c478a1",
  1770 => x"db03a9b7",
  1771 => x"48d4ff87",
  1772 => x"bfd8dec2",
  1773 => x"d4dec278",
  1774 => x"dec249bf",
  1775 => x"a1c148d4",
  1776 => x"b7c0c478",
  1777 => x"87e504a9",
  1778 => x"c848d0ff",
  1779 => x"e0dec278",
  1780 => x"2678c048",
  1781 => x"0000004f",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00005f5f",
  1785 => x"03030000",
  1786 => x"00030300",
  1787 => x"7f7f1400",
  1788 => x"147f7f14",
  1789 => x"2e240000",
  1790 => x"123a6b6b",
  1791 => x"366a4c00",
  1792 => x"32566c18",
  1793 => x"4f7e3000",
  1794 => x"683a7759",
  1795 => x"04000040",
  1796 => x"00000307",
  1797 => x"1c000000",
  1798 => x"0041633e",
  1799 => x"41000000",
  1800 => x"001c3e63",
  1801 => x"3e2a0800",
  1802 => x"2a3e1c1c",
  1803 => x"08080008",
  1804 => x"08083e3e",
  1805 => x"80000000",
  1806 => x"000060e0",
  1807 => x"08080000",
  1808 => x"08080808",
  1809 => x"00000000",
  1810 => x"00006060",
  1811 => x"30604000",
  1812 => x"03060c18",
  1813 => x"7f3e0001",
  1814 => x"3e7f4d59",
  1815 => x"06040000",
  1816 => x"00007f7f",
  1817 => x"63420000",
  1818 => x"464f5971",
  1819 => x"63220000",
  1820 => x"367f4949",
  1821 => x"161c1800",
  1822 => x"107f7f13",
  1823 => x"67270000",
  1824 => x"397d4545",
  1825 => x"7e3c0000",
  1826 => x"3079494b",
  1827 => x"01010000",
  1828 => x"070f7971",
  1829 => x"7f360000",
  1830 => x"367f4949",
  1831 => x"4f060000",
  1832 => x"1e3f6949",
  1833 => x"00000000",
  1834 => x"00006666",
  1835 => x"80000000",
  1836 => x"000066e6",
  1837 => x"08080000",
  1838 => x"22221414",
  1839 => x"14140000",
  1840 => x"14141414",
  1841 => x"22220000",
  1842 => x"08081414",
  1843 => x"03020000",
  1844 => x"060f5951",
  1845 => x"417f3e00",
  1846 => x"1e1f555d",
  1847 => x"7f7e0000",
  1848 => x"7e7f0909",
  1849 => x"7f7f0000",
  1850 => x"367f4949",
  1851 => x"3e1c0000",
  1852 => x"41414163",
  1853 => x"7f7f0000",
  1854 => x"1c3e6341",
  1855 => x"7f7f0000",
  1856 => x"41414949",
  1857 => x"7f7f0000",
  1858 => x"01010909",
  1859 => x"7f3e0000",
  1860 => x"7a7b4941",
  1861 => x"7f7f0000",
  1862 => x"7f7f0808",
  1863 => x"41000000",
  1864 => x"00417f7f",
  1865 => x"60200000",
  1866 => x"3f7f4040",
  1867 => x"087f7f00",
  1868 => x"4163361c",
  1869 => x"7f7f0000",
  1870 => x"40404040",
  1871 => x"067f7f00",
  1872 => x"7f7f060c",
  1873 => x"067f7f00",
  1874 => x"7f7f180c",
  1875 => x"7f3e0000",
  1876 => x"3e7f4141",
  1877 => x"7f7f0000",
  1878 => x"060f0909",
  1879 => x"417f3e00",
  1880 => x"407e7f61",
  1881 => x"7f7f0000",
  1882 => x"667f1909",
  1883 => x"6f260000",
  1884 => x"327b594d",
  1885 => x"01010000",
  1886 => x"01017f7f",
  1887 => x"7f3f0000",
  1888 => x"3f7f4040",
  1889 => x"3f0f0000",
  1890 => x"0f3f7070",
  1891 => x"307f7f00",
  1892 => x"7f7f3018",
  1893 => x"36634100",
  1894 => x"63361c1c",
  1895 => x"06030141",
  1896 => x"03067c7c",
  1897 => x"59716101",
  1898 => x"4143474d",
  1899 => x"7f000000",
  1900 => x"0041417f",
  1901 => x"06030100",
  1902 => x"6030180c",
  1903 => x"41000040",
  1904 => x"007f7f41",
  1905 => x"060c0800",
  1906 => x"080c0603",
  1907 => x"80808000",
  1908 => x"80808080",
  1909 => x"00000000",
  1910 => x"00040703",
  1911 => x"74200000",
  1912 => x"787c5454",
  1913 => x"7f7f0000",
  1914 => x"387c4444",
  1915 => x"7c380000",
  1916 => x"00444444",
  1917 => x"7c380000",
  1918 => x"7f7f4444",
  1919 => x"7c380000",
  1920 => x"185c5454",
  1921 => x"7e040000",
  1922 => x"0005057f",
  1923 => x"bc180000",
  1924 => x"7cfca4a4",
  1925 => x"7f7f0000",
  1926 => x"787c0404",
  1927 => x"00000000",
  1928 => x"00407d3d",
  1929 => x"80800000",
  1930 => x"007dfd80",
  1931 => x"7f7f0000",
  1932 => x"446c3810",
  1933 => x"00000000",
  1934 => x"00407f3f",
  1935 => x"0c7c7c00",
  1936 => x"787c0c18",
  1937 => x"7c7c0000",
  1938 => x"787c0404",
  1939 => x"7c380000",
  1940 => x"387c4444",
  1941 => x"fcfc0000",
  1942 => x"183c2424",
  1943 => x"3c180000",
  1944 => x"fcfc2424",
  1945 => x"7c7c0000",
  1946 => x"080c0404",
  1947 => x"5c480000",
  1948 => x"20745454",
  1949 => x"3f040000",
  1950 => x"0044447f",
  1951 => x"7c3c0000",
  1952 => x"7c7c4040",
  1953 => x"3c1c0000",
  1954 => x"1c3c6060",
  1955 => x"607c3c00",
  1956 => x"3c7c6030",
  1957 => x"386c4400",
  1958 => x"446c3810",
  1959 => x"bc1c0000",
  1960 => x"1c3c60e0",
  1961 => x"64440000",
  1962 => x"444c5c74",
  1963 => x"08080000",
  1964 => x"4141773e",
  1965 => x"00000000",
  1966 => x"00007f7f",
  1967 => x"41410000",
  1968 => x"08083e77",
  1969 => x"01010200",
  1970 => x"01020203",
  1971 => x"7f7f7f00",
  1972 => x"7f7f7f7f",
  1973 => x"1c080800",
  1974 => x"7f3e3e1c",
  1975 => x"3e7f7f7f",
  1976 => x"081c1c3e",
  1977 => x"18100008",
  1978 => x"10187c7c",
  1979 => x"30100000",
  1980 => x"10307c7c",
  1981 => x"60301000",
  1982 => x"061e7860",
  1983 => x"3c664200",
  1984 => x"42663c18",
  1985 => x"6a387800",
  1986 => x"386cc6c2",
  1987 => x"00006000",
  1988 => x"60000060",
  1989 => x"5b5e0e00",
  1990 => x"1e0e5d5c",
  1991 => x"dec24c71",
  1992 => x"c04dbfe5",
  1993 => x"741ec04b",
  1994 => x"87c702ab",
  1995 => x"c048a6c4",
  1996 => x"c487c578",
  1997 => x"78c148a6",
  1998 => x"731e66c4",
  1999 => x"87dfee49",
  2000 => x"e0c086c8",
  2001 => x"87eeef49",
  2002 => x"6a4aa5c4",
  2003 => x"87f0f049",
  2004 => x"cb87c6f1",
  2005 => x"c883c185",
  2006 => x"ff04abb7",
  2007 => x"262687c7",
  2008 => x"264c264d",
  2009 => x"1e4f264b",
  2010 => x"dec24a71",
  2011 => x"dec25ae9",
  2012 => x"78c748e9",
  2013 => x"87ddfe49",
  2014 => x"731e4f26",
  2015 => x"c04a711e",
  2016 => x"d303aab7",
  2017 => x"c3ccc287",
  2018 => x"87c405bf",
  2019 => x"87c24bc1",
  2020 => x"ccc24bc0",
  2021 => x"87c45bc7",
  2022 => x"5ac7ccc2",
  2023 => x"bfc3ccc2",
  2024 => x"c19ac14a",
  2025 => x"ec49a2c0",
  2026 => x"48fc87e8",
  2027 => x"bfc3ccc2",
  2028 => x"87effe78",
  2029 => x"c44a711e",
  2030 => x"49721e66",
  2031 => x"2687f9ea",
  2032 => x"ff1e4f26",
  2033 => x"ffc348d4",
  2034 => x"48d0ff78",
  2035 => x"ff78e1c0",
  2036 => x"78c148d4",
  2037 => x"30c44871",
  2038 => x"7808d4ff",
  2039 => x"c048d0ff",
  2040 => x"4f2678e0",
  2041 => x"5c5b5e0e",
  2042 => x"86f00e5d",
  2043 => x"c048a6c8",
  2044 => x"ec4b4d78",
  2045 => x"80fc7ebf",
  2046 => x"bfe5dec2",
  2047 => x"4cbfe878",
  2048 => x"bfc3ccc2",
  2049 => x"87cae349",
  2050 => x"cb49eecb",
  2051 => x"a6d087fd",
  2052 => x"e649c758",
  2053 => x"987087ff",
  2054 => x"6e87c805",
  2055 => x"0299c149",
  2056 => x"c187c3c1",
  2057 => x"7ebfec4b",
  2058 => x"bfc3ccc2",
  2059 => x"87e2e249",
  2060 => x"cb4966cc",
  2061 => x"987087e1",
  2062 => x"c287d802",
  2063 => x"49bffbcb",
  2064 => x"cbc2b9c1",
  2065 => x"fd7159ff",
  2066 => x"eecb87f8",
  2067 => x"87fbca49",
  2068 => x"c758a6d0",
  2069 => x"87fde549",
  2070 => x"ff059870",
  2071 => x"496e87c5",
  2072 => x"fe0599c1",
  2073 => x"9b7387fd",
  2074 => x"ff87d002",
  2075 => x"87cafc49",
  2076 => x"e549dac1",
  2077 => x"a6c887df",
  2078 => x"c278c148",
  2079 => x"05bfc3cc",
  2080 => x"c387e9c0",
  2081 => x"cce549fd",
  2082 => x"49fac387",
  2083 => x"7487c6e5",
  2084 => x"99ffc349",
  2085 => x"49c01e71",
  2086 => x"7487d9fc",
  2087 => x"29b7c849",
  2088 => x"49c11e71",
  2089 => x"c887cdfc",
  2090 => x"87f9c786",
  2091 => x"ffc34974",
  2092 => x"2cb7c899",
  2093 => x"9c74b471",
  2094 => x"c287dd02",
  2095 => x"49bfffcb",
  2096 => x"7087d4c9",
  2097 => x"87c40598",
  2098 => x"87d24cc0",
  2099 => x"c849e0c2",
  2100 => x"ccc287f9",
  2101 => x"87c658c3",
  2102 => x"48ffcbc2",
  2103 => x"497478c0",
  2104 => x"ce0599c2",
  2105 => x"49ebc387",
  2106 => x"7087eae3",
  2107 => x"0299c249",
  2108 => x"fb87c2c0",
  2109 => x"c149744d",
  2110 => x"87ce0599",
  2111 => x"e349f4c3",
  2112 => x"497087d3",
  2113 => x"c00299c2",
  2114 => x"4dfa87c2",
  2115 => x"99c84974",
  2116 => x"c387cd05",
  2117 => x"fce249f5",
  2118 => x"c2497087",
  2119 => x"87d90299",
  2120 => x"bfe9dec2",
  2121 => x"87cac002",
  2122 => x"c288c148",
  2123 => x"c058edde",
  2124 => x"4dff87c2",
  2125 => x"c148a6c8",
  2126 => x"c4497478",
  2127 => x"cdc00599",
  2128 => x"49f2c387",
  2129 => x"7087cee2",
  2130 => x"0299c249",
  2131 => x"dec287df",
  2132 => x"487ebfe9",
  2133 => x"03a8b7c7",
  2134 => x"6e87cbc0",
  2135 => x"c280c148",
  2136 => x"c058edde",
  2137 => x"4dfe87c2",
  2138 => x"c148a6c8",
  2139 => x"49fdc378",
  2140 => x"7087e2e1",
  2141 => x"0299c249",
  2142 => x"c287d8c0",
  2143 => x"02bfe9de",
  2144 => x"c287c9c0",
  2145 => x"c048e9de",
  2146 => x"87c2c078",
  2147 => x"a6c84dfd",
  2148 => x"c378c148",
  2149 => x"fce049fa",
  2150 => x"c2497087",
  2151 => x"dcc00299",
  2152 => x"e9dec287",
  2153 => x"b7c748bf",
  2154 => x"c9c003a8",
  2155 => x"e9dec287",
  2156 => x"c078c748",
  2157 => x"4dfc87c2",
  2158 => x"c148a6c8",
  2159 => x"adb7c078",
  2160 => x"87d0c003",
  2161 => x"c14a66c4",
  2162 => x"026a82d8",
  2163 => x"4b87c5c0",
  2164 => x"0f734975",
  2165 => x"dec24bc0",
  2166 => x"50c048e4",
  2167 => x"c449eecb",
  2168 => x"a6d087e9",
  2169 => x"e4dec258",
  2170 => x"c105bf97",
  2171 => x"497487de",
  2172 => x"0599f0c3",
  2173 => x"c187cdc0",
  2174 => x"dfff49da",
  2175 => x"987087d7",
  2176 => x"87c8c102",
  2177 => x"bfe84bc1",
  2178 => x"ffc3494c",
  2179 => x"2cb7c899",
  2180 => x"ccc2b471",
  2181 => x"ff49bfc3",
  2182 => x"cc87f7da",
  2183 => x"f6c34966",
  2184 => x"02987087",
  2185 => x"c287c6c0",
  2186 => x"c148e4de",
  2187 => x"e4dec250",
  2188 => x"c005bf97",
  2189 => x"497487d6",
  2190 => x"0599f0c3",
  2191 => x"c187c5ff",
  2192 => x"deff49da",
  2193 => x"987087cf",
  2194 => x"87f8fe05",
  2195 => x"c0029b73",
  2196 => x"a6cc87e0",
  2197 => x"e9dec248",
  2198 => x"66cc78bf",
  2199 => x"c491cb49",
  2200 => x"80714866",
  2201 => x"bf6e7e70",
  2202 => x"87c6c002",
  2203 => x"4966cc4b",
  2204 => x"66c80f73",
  2205 => x"87c8c002",
  2206 => x"bfe9dec2",
  2207 => x"87d5f249",
  2208 => x"bfc7ccc2",
  2209 => x"87ddc002",
  2210 => x"87cbc249",
  2211 => x"c0029870",
  2212 => x"dec287d3",
  2213 => x"f149bfe9",
  2214 => x"49c087fb",
  2215 => x"c287dbf3",
  2216 => x"c048c7cc",
  2217 => x"f28ef078",
  2218 => x"5e0e87f5",
  2219 => x"0e5d5c5b",
  2220 => x"c24c711e",
  2221 => x"49bfe5de",
  2222 => x"4da1cdc1",
  2223 => x"6981d1c1",
  2224 => x"029c747e",
  2225 => x"a5c487cf",
  2226 => x"c27b744b",
  2227 => x"49bfe5de",
  2228 => x"6e87d4f2",
  2229 => x"059c747b",
  2230 => x"4bc087c4",
  2231 => x"4bc187c2",
  2232 => x"d5f24973",
  2233 => x"0266d487",
  2234 => x"de4987c7",
  2235 => x"c24a7087",
  2236 => x"c24ac087",
  2237 => x"265acbcc",
  2238 => x"0087e4f1",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"1e000000",
  2243 => x"c8ff4a71",
  2244 => x"a17249bf",
  2245 => x"1e4f2648",
  2246 => x"89bfc8ff",
  2247 => x"c0c0c0fe",
  2248 => x"01a9c0c0",
  2249 => x"4ac087c4",
  2250 => x"4ac187c2",
  2251 => x"4f264872",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
