library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e8dec287",
    12 => x"86c0c84e",
    13 => x"49e8dec2",
    14 => x"48e8ccc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c6dc",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c348724c",
    72 => x"7c7098ff",
    73 => x"bfe8ccc2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"ffc34871",
    79 => x"d07c7098",
    80 => x"29d04966",
    81 => x"ffc34871",
    82 => x"d07c7098",
    83 => x"29c84966",
    84 => x"ffc34871",
    85 => x"d07c7098",
    86 => x"ffc34866",
    87 => x"727c7098",
    88 => x"7129d049",
    89 => x"98ffc348",
    90 => x"4b6c7c70",
    91 => x"4dfff0c9",
    92 => x"05abffc3",
    93 => x"ffc387d0",
    94 => x"c14b6c7c",
    95 => x"87c6028d",
    96 => x"02abffc3",
    97 => x"487387f0",
    98 => x"1e87fffd",
    99 => x"d4ff49c0",
   100 => x"78ffc348",
   101 => x"c8c381c1",
   102 => x"f104a9b7",
   103 => x"1e4f2687",
   104 => x"87e71e73",
   105 => x"4bdff8c4",
   106 => x"ffc01ec0",
   107 => x"49f7c1f0",
   108 => x"c487dffd",
   109 => x"05a8c186",
   110 => x"ff87eac0",
   111 => x"ffc348d4",
   112 => x"c0c0c178",
   113 => x"1ec0c0c0",
   114 => x"c1f0e1c0",
   115 => x"c1fd49e9",
   116 => x"7086c487",
   117 => x"87ca0598",
   118 => x"c348d4ff",
   119 => x"48c178ff",
   120 => x"e6fe87cb",
   121 => x"058bc187",
   122 => x"c087fdfe",
   123 => x"87defc48",
   124 => x"ff1e731e",
   125 => x"ffc348d4",
   126 => x"c04bd378",
   127 => x"f0ffc01e",
   128 => x"fc49c1c1",
   129 => x"86c487cc",
   130 => x"ca059870",
   131 => x"48d4ff87",
   132 => x"c178ffc3",
   133 => x"fd87cb48",
   134 => x"8bc187f1",
   135 => x"87dbff05",
   136 => x"e9fb48c0",
   137 => x"5b5e0e87",
   138 => x"d4ff0e5c",
   139 => x"87dbfd4c",
   140 => x"c01eeac6",
   141 => x"c8c1f0e1",
   142 => x"87d6fb49",
   143 => x"a8c186c4",
   144 => x"fe87c802",
   145 => x"48c087ea",
   146 => x"fa87e2c1",
   147 => x"497087d2",
   148 => x"99ffffcf",
   149 => x"02a9eac6",
   150 => x"d3fe87c8",
   151 => x"c148c087",
   152 => x"ffc387cb",
   153 => x"4bf1c07c",
   154 => x"7087f4fc",
   155 => x"ebc00298",
   156 => x"c01ec087",
   157 => x"fac1f0ff",
   158 => x"87d6fa49",
   159 => x"987086c4",
   160 => x"c387d905",
   161 => x"496c7cff",
   162 => x"7c7cffc3",
   163 => x"c0c17c7c",
   164 => x"87c40299",
   165 => x"87d548c1",
   166 => x"87d148c0",
   167 => x"c405abc2",
   168 => x"c848c087",
   169 => x"058bc187",
   170 => x"c087fdfe",
   171 => x"87dcf948",
   172 => x"c21e731e",
   173 => x"c148e8cc",
   174 => x"ff4bc778",
   175 => x"78c248d0",
   176 => x"ff87c8fb",
   177 => x"78c348d0",
   178 => x"e5c01ec0",
   179 => x"49c0c1d0",
   180 => x"c487fff8",
   181 => x"05a8c186",
   182 => x"c24b87c1",
   183 => x"87c505ab",
   184 => x"f9c048c0",
   185 => x"058bc187",
   186 => x"fc87d0ff",
   187 => x"ccc287f7",
   188 => x"987058ec",
   189 => x"c187cd05",
   190 => x"f0ffc01e",
   191 => x"f849d0c1",
   192 => x"86c487d0",
   193 => x"c348d4ff",
   194 => x"fdc278ff",
   195 => x"f0ccc287",
   196 => x"48d0ff58",
   197 => x"d4ff78c2",
   198 => x"78ffc348",
   199 => x"edf748c1",
   200 => x"5b5e0e87",
   201 => x"710e5d5c",
   202 => x"c54cc04b",
   203 => x"4adfcdee",
   204 => x"c348d4ff",
   205 => x"486878ff",
   206 => x"05a8fec3",
   207 => x"ff87fec0",
   208 => x"9b734dd4",
   209 => x"d087cc02",
   210 => x"49731e66",
   211 => x"c487e8f5",
   212 => x"ff87d686",
   213 => x"d1c448d0",
   214 => x"7dffc378",
   215 => x"c14866d0",
   216 => x"58a6d488",
   217 => x"f0059870",
   218 => x"48d4ff87",
   219 => x"7878ffc3",
   220 => x"c5059b73",
   221 => x"48d0ff87",
   222 => x"4ac178d0",
   223 => x"058ac14c",
   224 => x"7487edfe",
   225 => x"87c2f648",
   226 => x"711e731e",
   227 => x"ff4bc04a",
   228 => x"ffc348d4",
   229 => x"48d0ff78",
   230 => x"ff78c3c4",
   231 => x"ffc348d4",
   232 => x"c01e7278",
   233 => x"d1c1f0ff",
   234 => x"87e6f549",
   235 => x"987086c4",
   236 => x"c887d205",
   237 => x"66cc1ec0",
   238 => x"87e5fd49",
   239 => x"4b7086c4",
   240 => x"c248d0ff",
   241 => x"f5487378",
   242 => x"5e0e87c4",
   243 => x"0e5d5c5b",
   244 => x"ffc01ec0",
   245 => x"49c9c1f0",
   246 => x"d287f7f4",
   247 => x"f0ccc21e",
   248 => x"87fdfc49",
   249 => x"4cc086c8",
   250 => x"b7d284c1",
   251 => x"87f804ac",
   252 => x"97f0ccc2",
   253 => x"c0c349bf",
   254 => x"a9c0c199",
   255 => x"87e7c005",
   256 => x"97f7ccc2",
   257 => x"31d049bf",
   258 => x"97f8ccc2",
   259 => x"32c84abf",
   260 => x"ccc2b172",
   261 => x"4abf97f9",
   262 => x"cf4c71b1",
   263 => x"9cffffff",
   264 => x"34ca84c1",
   265 => x"c287e7c1",
   266 => x"bf97f9cc",
   267 => x"c631c149",
   268 => x"faccc299",
   269 => x"c74abf97",
   270 => x"b1722ab7",
   271 => x"97f5ccc2",
   272 => x"cf4d4abf",
   273 => x"f6ccc29d",
   274 => x"c34abf97",
   275 => x"c232ca9a",
   276 => x"bf97f7cc",
   277 => x"7333c24b",
   278 => x"f8ccc2b2",
   279 => x"c34bbf97",
   280 => x"b7c69bc0",
   281 => x"c2b2732b",
   282 => x"7148c181",
   283 => x"c1497030",
   284 => x"70307548",
   285 => x"c14c724d",
   286 => x"c8947184",
   287 => x"06adb7c0",
   288 => x"34c187cc",
   289 => x"c0c82db7",
   290 => x"ff01adb7",
   291 => x"487487f4",
   292 => x"0e87f7f1",
   293 => x"5d5c5b5e",
   294 => x"c286f80e",
   295 => x"c048d6d5",
   296 => x"cecdc278",
   297 => x"fb49c01e",
   298 => x"86c487de",
   299 => x"c5059870",
   300 => x"c948c087",
   301 => x"4dc087c0",
   302 => x"edc07ec1",
   303 => x"c249bfe6",
   304 => x"714ac4ce",
   305 => x"e0ee4bc8",
   306 => x"05987087",
   307 => x"7ec087c2",
   308 => x"bfe2edc0",
   309 => x"e0cec249",
   310 => x"4bc8714a",
   311 => x"7087caee",
   312 => x"87c20598",
   313 => x"026e7ec0",
   314 => x"c287fdc0",
   315 => x"4dbfd4d4",
   316 => x"9fccd5c2",
   317 => x"c5487ebf",
   318 => x"05a8ead6",
   319 => x"d4c287c7",
   320 => x"ce4dbfd4",
   321 => x"ca486e87",
   322 => x"02a8d5e9",
   323 => x"48c087c5",
   324 => x"c287e3c7",
   325 => x"751ececd",
   326 => x"87ecf949",
   327 => x"987086c4",
   328 => x"c087c505",
   329 => x"87cec748",
   330 => x"bfe2edc0",
   331 => x"e0cec249",
   332 => x"4bc8714a",
   333 => x"7087f2ec",
   334 => x"87c80598",
   335 => x"48d6d5c2",
   336 => x"87da78c1",
   337 => x"bfe6edc0",
   338 => x"c4cec249",
   339 => x"4bc8714a",
   340 => x"7087d6ec",
   341 => x"c5c00298",
   342 => x"c648c087",
   343 => x"d5c287d8",
   344 => x"49bf97cc",
   345 => x"05a9d5c1",
   346 => x"c287cdc0",
   347 => x"bf97cdd5",
   348 => x"a9eac249",
   349 => x"87c5c002",
   350 => x"f9c548c0",
   351 => x"cecdc287",
   352 => x"487ebf97",
   353 => x"02a8e9c3",
   354 => x"6e87cec0",
   355 => x"a8ebc348",
   356 => x"87c5c002",
   357 => x"ddc548c0",
   358 => x"d9cdc287",
   359 => x"9949bf97",
   360 => x"87ccc005",
   361 => x"97dacdc2",
   362 => x"a9c249bf",
   363 => x"87c5c002",
   364 => x"c1c548c0",
   365 => x"dbcdc287",
   366 => x"c248bf97",
   367 => x"7058d2d5",
   368 => x"88c1484c",
   369 => x"58d6d5c2",
   370 => x"97dccdc2",
   371 => x"817549bf",
   372 => x"97ddcdc2",
   373 => x"32c84abf",
   374 => x"c27ea172",
   375 => x"6e48e3d9",
   376 => x"decdc278",
   377 => x"c848bf97",
   378 => x"d5c258a6",
   379 => x"c202bfd6",
   380 => x"edc087cf",
   381 => x"c249bfe2",
   382 => x"714ae0ce",
   383 => x"e8e94bc8",
   384 => x"02987087",
   385 => x"c087c5c0",
   386 => x"87eac348",
   387 => x"bfced5c2",
   388 => x"f7d9c24c",
   389 => x"f3cdc25c",
   390 => x"c849bf97",
   391 => x"f2cdc231",
   392 => x"a14abf97",
   393 => x"f4cdc249",
   394 => x"d04abf97",
   395 => x"49a17232",
   396 => x"97f5cdc2",
   397 => x"32d84abf",
   398 => x"c449a172",
   399 => x"d9c29166",
   400 => x"c281bfe3",
   401 => x"c259ebd9",
   402 => x"bf97fbcd",
   403 => x"c232c84a",
   404 => x"bf97facd",
   405 => x"c24aa24b",
   406 => x"bf97fccd",
   407 => x"7333d04b",
   408 => x"cdc24aa2",
   409 => x"4bbf97fd",
   410 => x"33d89bcf",
   411 => x"c24aa273",
   412 => x"c25aefd9",
   413 => x"c292748a",
   414 => x"7248efd9",
   415 => x"c1c178a1",
   416 => x"e0cdc287",
   417 => x"c849bf97",
   418 => x"dfcdc231",
   419 => x"a14abf97",
   420 => x"c731c549",
   421 => x"29c981ff",
   422 => x"59f7d9c2",
   423 => x"97e5cdc2",
   424 => x"32c84abf",
   425 => x"97e4cdc2",
   426 => x"4aa24bbf",
   427 => x"6e9266c4",
   428 => x"f3d9c282",
   429 => x"ebd9c25a",
   430 => x"c278c048",
   431 => x"7248e7d9",
   432 => x"d9c278a1",
   433 => x"d9c248f7",
   434 => x"c278bfeb",
   435 => x"c248fbd9",
   436 => x"78bfefd9",
   437 => x"bfd6d5c2",
   438 => x"87c9c002",
   439 => x"30c44874",
   440 => x"c9c07e70",
   441 => x"f3d9c287",
   442 => x"30c448bf",
   443 => x"d5c27e70",
   444 => x"786e48da",
   445 => x"8ef848c1",
   446 => x"4c264d26",
   447 => x"4f264b26",
   448 => x"5c5b5e0e",
   449 => x"4a710e5d",
   450 => x"bfd6d5c2",
   451 => x"7287cb02",
   452 => x"722bc74b",
   453 => x"9dffc14d",
   454 => x"4b7287c9",
   455 => x"4d722bc8",
   456 => x"c29dffc3",
   457 => x"83bfe3d9",
   458 => x"bfdeedc0",
   459 => x"87d902ab",
   460 => x"5be2edc0",
   461 => x"1ececdc2",
   462 => x"cbf14973",
   463 => x"7086c487",
   464 => x"87c50598",
   465 => x"e6c048c0",
   466 => x"d6d5c287",
   467 => x"87d202bf",
   468 => x"91c44975",
   469 => x"81cecdc2",
   470 => x"ffcf4c69",
   471 => x"9cffffff",
   472 => x"497587cb",
   473 => x"cdc291c2",
   474 => x"699f81ce",
   475 => x"fe48744c",
   476 => x"5e0e87c6",
   477 => x"0e5d5c5b",
   478 => x"4c7186f8",
   479 => x"87c5059c",
   480 => x"c0c348c0",
   481 => x"7ea4c887",
   482 => x"d878c048",
   483 => x"87c70266",
   484 => x"bf9766d8",
   485 => x"c087c505",
   486 => x"87e9c248",
   487 => x"49c11ec0",
   488 => x"87e3c749",
   489 => x"4d7086c4",
   490 => x"c2c1029d",
   491 => x"ded5c287",
   492 => x"4966d84a",
   493 => x"7087d7e2",
   494 => x"f2c00298",
   495 => x"d84a7587",
   496 => x"4bcb4966",
   497 => x"7087fce2",
   498 => x"e2c00298",
   499 => x"751ec087",
   500 => x"87c7029d",
   501 => x"c048a6c8",
   502 => x"c887c578",
   503 => x"78c148a6",
   504 => x"c64966c8",
   505 => x"86c487e1",
   506 => x"059d4d70",
   507 => x"7587fefe",
   508 => x"cec1029d",
   509 => x"49a5dc87",
   510 => x"7869486e",
   511 => x"c449a5da",
   512 => x"a4c448a6",
   513 => x"48699f78",
   514 => x"780866c4",
   515 => x"bfd6d5c2",
   516 => x"d487d202",
   517 => x"699f49a5",
   518 => x"ffffc049",
   519 => x"d0487199",
   520 => x"c27e7030",
   521 => x"6e7ec087",
   522 => x"bf66c448",
   523 => x"0866c480",
   524 => x"cc7cc078",
   525 => x"66c449a4",
   526 => x"a4d079bf",
   527 => x"c179c049",
   528 => x"c087c248",
   529 => x"fa8ef848",
   530 => x"5e0e87ee",
   531 => x"710e5c5b",
   532 => x"c1029c4c",
   533 => x"a4c887cb",
   534 => x"c1026949",
   535 => x"496c87c3",
   536 => x"714866cc",
   537 => x"58a6d080",
   538 => x"d5c2b970",
   539 => x"ff4abfd2",
   540 => x"719972ba",
   541 => x"e5c00299",
   542 => x"4ba4c487",
   543 => x"fff9496b",
   544 => x"c27b7087",
   545 => x"49bfced5",
   546 => x"7c71816c",
   547 => x"c2b966cc",
   548 => x"4abfd2d5",
   549 => x"9972baff",
   550 => x"ff059971",
   551 => x"66cc87db",
   552 => x"87d6f97c",
   553 => x"711e731e",
   554 => x"c7029b4b",
   555 => x"49a3c887",
   556 => x"87c50569",
   557 => x"f6c048c0",
   558 => x"e7d9c287",
   559 => x"a3c449bf",
   560 => x"c24a6a4a",
   561 => x"ced5c28a",
   562 => x"a17292bf",
   563 => x"d2d5c249",
   564 => x"9a6b4abf",
   565 => x"c049a172",
   566 => x"c859e2ed",
   567 => x"ea711e66",
   568 => x"86c487e6",
   569 => x"c4059870",
   570 => x"c248c087",
   571 => x"f848c187",
   572 => x"731e87ca",
   573 => x"9b4b711e",
   574 => x"87e4c002",
   575 => x"5bfbd9c2",
   576 => x"8ac24a73",
   577 => x"bfced5c2",
   578 => x"d9c29249",
   579 => x"7248bfe7",
   580 => x"ffd9c280",
   581 => x"c4487158",
   582 => x"ded5c230",
   583 => x"87edc058",
   584 => x"48f7d9c2",
   585 => x"bfebd9c2",
   586 => x"fbd9c278",
   587 => x"efd9c248",
   588 => x"d5c278bf",
   589 => x"c902bfd6",
   590 => x"ced5c287",
   591 => x"31c449bf",
   592 => x"d9c287c7",
   593 => x"c449bff3",
   594 => x"ded5c231",
   595 => x"87ecf659",
   596 => x"5c5b5e0e",
   597 => x"c04a710e",
   598 => x"029a724b",
   599 => x"da87e0c0",
   600 => x"699f49a2",
   601 => x"d6d5c24b",
   602 => x"87cf02bf",
   603 => x"9f49a2d4",
   604 => x"c04c4969",
   605 => x"d09cffff",
   606 => x"c087c234",
   607 => x"73b3744c",
   608 => x"87eefd49",
   609 => x"0e87f3f5",
   610 => x"5d5c5b5e",
   611 => x"7186f40e",
   612 => x"727ec04a",
   613 => x"87d8029a",
   614 => x"48cacdc2",
   615 => x"cdc278c0",
   616 => x"d9c248c2",
   617 => x"c278bffb",
   618 => x"c248c6cd",
   619 => x"78bff7d9",
   620 => x"48ebd5c2",
   621 => x"d5c250c0",
   622 => x"c249bfda",
   623 => x"4abfcacd",
   624 => x"c403aa71",
   625 => x"497287c9",
   626 => x"c00599cf",
   627 => x"edc087e9",
   628 => x"cdc248de",
   629 => x"c278bfc2",
   630 => x"c21ececd",
   631 => x"49bfc2cd",
   632 => x"48c2cdc2",
   633 => x"7178a1c1",
   634 => x"c487dde6",
   635 => x"daedc086",
   636 => x"cecdc248",
   637 => x"c087cc78",
   638 => x"48bfdaed",
   639 => x"c080e0c0",
   640 => x"c258deed",
   641 => x"48bfcacd",
   642 => x"cdc280c1",
   643 => x"5a2758ce",
   644 => x"bf00000b",
   645 => x"9d4dbf97",
   646 => x"87e3c202",
   647 => x"02ade5c3",
   648 => x"c087dcc2",
   649 => x"4bbfdaed",
   650 => x"1149a3cb",
   651 => x"05accf4c",
   652 => x"7587d2c1",
   653 => x"c199df49",
   654 => x"c291cd89",
   655 => x"c181ded5",
   656 => x"51124aa3",
   657 => x"124aa3c3",
   658 => x"4aa3c551",
   659 => x"a3c75112",
   660 => x"c951124a",
   661 => x"51124aa3",
   662 => x"124aa3ce",
   663 => x"4aa3d051",
   664 => x"a3d25112",
   665 => x"d451124a",
   666 => x"51124aa3",
   667 => x"124aa3d6",
   668 => x"4aa3d851",
   669 => x"a3dc5112",
   670 => x"de51124a",
   671 => x"51124aa3",
   672 => x"fac07ec1",
   673 => x"c8497487",
   674 => x"ebc00599",
   675 => x"d0497487",
   676 => x"87d10599",
   677 => x"c00266dc",
   678 => x"497387cb",
   679 => x"700f66dc",
   680 => x"d3c00298",
   681 => x"c0056e87",
   682 => x"d5c287c6",
   683 => x"50c048de",
   684 => x"bfdaedc0",
   685 => x"87ddc248",
   686 => x"48ebd5c2",
   687 => x"c27e50c0",
   688 => x"49bfdad5",
   689 => x"bfcacdc2",
   690 => x"04aa714a",
   691 => x"c287f7fb",
   692 => x"05bffbd9",
   693 => x"c287c8c0",
   694 => x"02bfd6d5",
   695 => x"c287f4c1",
   696 => x"49bfc6cd",
   697 => x"c287d9f0",
   698 => x"c458cacd",
   699 => x"cdc248a6",
   700 => x"c278bfc6",
   701 => x"02bfd6d5",
   702 => x"c487d8c0",
   703 => x"ffcf4966",
   704 => x"99f8ffff",
   705 => x"c5c002a9",
   706 => x"c04cc087",
   707 => x"4cc187e1",
   708 => x"c487dcc0",
   709 => x"ffcf4966",
   710 => x"02a999f8",
   711 => x"c887c8c0",
   712 => x"78c048a6",
   713 => x"c887c5c0",
   714 => x"78c148a6",
   715 => x"744c66c8",
   716 => x"dec0059c",
   717 => x"4966c487",
   718 => x"d5c289c2",
   719 => x"c291bfce",
   720 => x"48bfe7d9",
   721 => x"cdc28071",
   722 => x"cdc258c6",
   723 => x"78c048ca",
   724 => x"c087e3f9",
   725 => x"ee8ef448",
   726 => x"000087de",
   727 => x"ffff0000",
   728 => x"0b6affff",
   729 => x"0b730000",
   730 => x"41460000",
   731 => x"20323354",
   732 => x"46002020",
   733 => x"36315441",
   734 => x"00202020",
   735 => x"48d4ff1e",
   736 => x"6878ffc3",
   737 => x"1e4f2648",
   738 => x"c348d4ff",
   739 => x"d0ff78ff",
   740 => x"78e1c048",
   741 => x"d448d4ff",
   742 => x"ffd9c278",
   743 => x"bfd4ff48",
   744 => x"1e4f2650",
   745 => x"c048d0ff",
   746 => x"4f2678e0",
   747 => x"87ccff1e",
   748 => x"02994970",
   749 => x"fbc087c6",
   750 => x"87f105a9",
   751 => x"4f264871",
   752 => x"5c5b5e0e",
   753 => x"c04b710e",
   754 => x"87f0fe4c",
   755 => x"02994970",
   756 => x"c087f9c0",
   757 => x"c002a9ec",
   758 => x"fbc087f2",
   759 => x"ebc002a9",
   760 => x"b766cc87",
   761 => x"87c703ac",
   762 => x"c20266d0",
   763 => x"71537187",
   764 => x"87c20299",
   765 => x"c3fe84c1",
   766 => x"99497087",
   767 => x"c087cd02",
   768 => x"c702a9ec",
   769 => x"a9fbc087",
   770 => x"87d5ff05",
   771 => x"c30266d0",
   772 => x"7b97c087",
   773 => x"05a9ecc0",
   774 => x"4a7487c4",
   775 => x"4a7487c5",
   776 => x"728a0ac0",
   777 => x"2687c248",
   778 => x"264c264d",
   779 => x"1e4f264b",
   780 => x"7087c9fd",
   781 => x"a9f0c049",
   782 => x"c087c904",
   783 => x"c301a9f9",
   784 => x"89f0c087",
   785 => x"04a9c1c1",
   786 => x"dac187c9",
   787 => x"87c301a9",
   788 => x"7189f7c0",
   789 => x"0e4f2648",
   790 => x"5d5c5b5e",
   791 => x"7186f80e",
   792 => x"fc4dc04c",
   793 => x"4bc087e1",
   794 => x"97f6f3c0",
   795 => x"a9c049bf",
   796 => x"fc87cf04",
   797 => x"83c187f6",
   798 => x"97f6f3c0",
   799 => x"06ab49bf",
   800 => x"f3c087f1",
   801 => x"02bf97f6",
   802 => x"effb87cf",
   803 => x"99497087",
   804 => x"c087c602",
   805 => x"f105a9ec",
   806 => x"fb4bc087",
   807 => x"7e7087de",
   808 => x"c887d9fb",
   809 => x"d3fb58a6",
   810 => x"c14a7087",
   811 => x"49a4c883",
   812 => x"6e496997",
   813 => x"87da05a9",
   814 => x"9749a4c9",
   815 => x"66c44969",
   816 => x"87ce05a9",
   817 => x"9749a4ca",
   818 => x"05aa4969",
   819 => x"4dc187c4",
   820 => x"486e87d4",
   821 => x"02a8ecc0",
   822 => x"486e87c8",
   823 => x"05a8fbc0",
   824 => x"4bc087c4",
   825 => x"9d754dc1",
   826 => x"87effe02",
   827 => x"7387f4fa",
   828 => x"fc8ef848",
   829 => x"0e0087f1",
   830 => x"5d5c5b5e",
   831 => x"7186f80e",
   832 => x"4bd4ff7e",
   833 => x"dac21e6e",
   834 => x"e5e949c4",
   835 => x"7086c487",
   836 => x"eac40298",
   837 => x"ddddc187",
   838 => x"496e4dbf",
   839 => x"c887f8fc",
   840 => x"987058a6",
   841 => x"c487c505",
   842 => x"78c148a6",
   843 => x"c548d0ff",
   844 => x"7bd5c178",
   845 => x"c14966c4",
   846 => x"c131c689",
   847 => x"bf97dbdd",
   848 => x"b071484a",
   849 => x"d0ff7b70",
   850 => x"c278c448",
   851 => x"bf97ffd9",
   852 => x"0299d049",
   853 => x"78c587d7",
   854 => x"c07bd6c1",
   855 => x"7bffc34a",
   856 => x"e0c082c1",
   857 => x"87f504aa",
   858 => x"c448d0ff",
   859 => x"7bffc378",
   860 => x"c548d0ff",
   861 => x"7bd3c178",
   862 => x"78c47bc1",
   863 => x"06adb7c0",
   864 => x"c287ebc2",
   865 => x"4cbfccda",
   866 => x"c2029c8d",
   867 => x"cdc287c2",
   868 => x"a6c47ece",
   869 => x"78c0c848",
   870 => x"acb7c08c",
   871 => x"c887c603",
   872 => x"c078a4c0",
   873 => x"ffd9c24c",
   874 => x"d049bf97",
   875 => x"87d00299",
   876 => x"dac21ec0",
   877 => x"ebeb49c4",
   878 => x"7086c487",
   879 => x"87f5c04a",
   880 => x"1ececdc2",
   881 => x"49c4dac2",
   882 => x"c487d9eb",
   883 => x"ff4a7086",
   884 => x"c5c848d0",
   885 => x"7bd4c178",
   886 => x"7bbf976e",
   887 => x"80c1486e",
   888 => x"66c47e70",
   889 => x"c888c148",
   890 => x"987058a6",
   891 => x"87e8ff05",
   892 => x"c448d0ff",
   893 => x"059a7278",
   894 => x"48c087c5",
   895 => x"c187c2c1",
   896 => x"c4dac21e",
   897 => x"87c2e949",
   898 => x"9c7486c4",
   899 => x"87fefd05",
   900 => x"06adb7c0",
   901 => x"dac287d1",
   902 => x"78c048c4",
   903 => x"78c080d0",
   904 => x"dac280f4",
   905 => x"c078bfd0",
   906 => x"fd01adb7",
   907 => x"d0ff87d5",
   908 => x"c178c548",
   909 => x"7bc07bd3",
   910 => x"48c178c4",
   911 => x"c087c2c0",
   912 => x"268ef848",
   913 => x"264c264d",
   914 => x"0e4f264b",
   915 => x"5d5c5b5e",
   916 => x"4b711e0e",
   917 => x"ab4d4cc0",
   918 => x"87e8c004",
   919 => x"1ed7f1c0",
   920 => x"c4029d75",
   921 => x"c24ac087",
   922 => x"724ac187",
   923 => x"87d7ec49",
   924 => x"7e7086c4",
   925 => x"056e84c1",
   926 => x"4c7387c2",
   927 => x"ac7385c1",
   928 => x"87d8ff06",
   929 => x"fe26486e",
   930 => x"711e87f9",
   931 => x"0566c44a",
   932 => x"497287c5",
   933 => x"2687e0f9",
   934 => x"5b5e0e4f",
   935 => x"1e0e5d5c",
   936 => x"de494c71",
   937 => x"ecdac291",
   938 => x"9785714d",
   939 => x"dcc1026d",
   940 => x"d8dac287",
   941 => x"817449bf",
   942 => x"87cffe71",
   943 => x"98487e70",
   944 => x"87f2c002",
   945 => x"4be0dac2",
   946 => x"49cb4a70",
   947 => x"87d7c7ff",
   948 => x"93cb4b74",
   949 => x"83efddc1",
   950 => x"fcc083c4",
   951 => x"49747bd1",
   952 => x"87e9c0c1",
   953 => x"ddc17b75",
   954 => x"49bf97dc",
   955 => x"e0dac21e",
   956 => x"87d6fe49",
   957 => x"497486c4",
   958 => x"87d1c0c1",
   959 => x"c1c149c0",
   960 => x"dac287f0",
   961 => x"78c048c0",
   962 => x"f9dd49c1",
   963 => x"f2fc2687",
   964 => x"616f4c87",
   965 => x"676e6964",
   966 => x"002e2e2e",
   967 => x"711e731e",
   968 => x"dac2494a",
   969 => x"7181bfd8",
   970 => x"7087e0fc",
   971 => x"c4029b4b",
   972 => x"dbe84987",
   973 => x"d8dac287",
   974 => x"c178c048",
   975 => x"87c6dd49",
   976 => x"1e87c4fc",
   977 => x"c0c149c0",
   978 => x"4f2687e8",
   979 => x"494a711e",
   980 => x"ddc191cb",
   981 => x"81c881ef",
   982 => x"dac24811",
   983 => x"dac258c4",
   984 => x"78c048d8",
   985 => x"dddc49c1",
   986 => x"1e4f2687",
   987 => x"d2029971",
   988 => x"c4dfc187",
   989 => x"f750c048",
   990 => x"ccfdc080",
   991 => x"e8ddc140",
   992 => x"c187ce78",
   993 => x"c148c0df",
   994 => x"fc78e1dd",
   995 => x"c3fdc080",
   996 => x"0e4f2678",
   997 => x"5d5c5b5e",
   998 => x"c286f40e",
   999 => x"c04dcecd",
  1000 => x"48a6c44c",
  1001 => x"dac278c0",
  1002 => x"c048bfd8",
  1003 => x"c0c106a8",
  1004 => x"cecdc287",
  1005 => x"c0029848",
  1006 => x"f1c087f7",
  1007 => x"66c81ed7",
  1008 => x"c487c702",
  1009 => x"78c048a6",
  1010 => x"a6c487c5",
  1011 => x"c478c148",
  1012 => x"f2e64966",
  1013 => x"7086c487",
  1014 => x"c484c14d",
  1015 => x"80c14866",
  1016 => x"c258a6c8",
  1017 => x"acbfd8da",
  1018 => x"7587c603",
  1019 => x"c9ff059d",
  1020 => x"754cc087",
  1021 => x"dcc3029d",
  1022 => x"d7f1c087",
  1023 => x"0266c81e",
  1024 => x"a6cc87c7",
  1025 => x"c578c048",
  1026 => x"48a6cc87",
  1027 => x"66cc78c1",
  1028 => x"87f3e549",
  1029 => x"7e7086c4",
  1030 => x"c2029848",
  1031 => x"cb4987e4",
  1032 => x"49699781",
  1033 => x"c10299d0",
  1034 => x"497487d4",
  1035 => x"ddc191cb",
  1036 => x"fcc081ef",
  1037 => x"81c879dc",
  1038 => x"7451ffc3",
  1039 => x"c291de49",
  1040 => x"714decda",
  1041 => x"97c1c285",
  1042 => x"49a5c17d",
  1043 => x"c251e0c0",
  1044 => x"bf97ded5",
  1045 => x"c187d202",
  1046 => x"4ba5c284",
  1047 => x"4aded5c2",
  1048 => x"c1ff49db",
  1049 => x"d9c187c1",
  1050 => x"49a5cd87",
  1051 => x"84c151c0",
  1052 => x"6e4ba5c2",
  1053 => x"ff49cb4a",
  1054 => x"c187ecc0",
  1055 => x"497487c4",
  1056 => x"ddc191cb",
  1057 => x"fac081ef",
  1058 => x"d5c279d9",
  1059 => x"02bf97de",
  1060 => x"497487d8",
  1061 => x"84c191de",
  1062 => x"4becdac2",
  1063 => x"d5c28371",
  1064 => x"49dd4ade",
  1065 => x"87fffffe",
  1066 => x"4b7487d8",
  1067 => x"dac293de",
  1068 => x"a3cb83ec",
  1069 => x"c151c049",
  1070 => x"4a6e7384",
  1071 => x"fffe49cb",
  1072 => x"66c487e5",
  1073 => x"c880c148",
  1074 => x"acc758a6",
  1075 => x"87c5c003",
  1076 => x"e4fc056e",
  1077 => x"f4487487",
  1078 => x"87e7f58e",
  1079 => x"711e731e",
  1080 => x"91cb494b",
  1081 => x"81efddc1",
  1082 => x"c14aa1c8",
  1083 => x"1248dbdd",
  1084 => x"4aa1c950",
  1085 => x"48f6f3c0",
  1086 => x"81ca5012",
  1087 => x"48dcddc1",
  1088 => x"ddc15011",
  1089 => x"49bf97dc",
  1090 => x"f549c01e",
  1091 => x"dac287fc",
  1092 => x"78de48c0",
  1093 => x"edd549c1",
  1094 => x"eaf42687",
  1095 => x"5b5e0e87",
  1096 => x"f40e5d5c",
  1097 => x"494d7186",
  1098 => x"ddc191cb",
  1099 => x"a1c881ef",
  1100 => x"7ea1ca4a",
  1101 => x"c248a6c4",
  1102 => x"78bfc8de",
  1103 => x"4bbf976e",
  1104 => x"734c66c4",
  1105 => x"cc48122c",
  1106 => x"9c7058a6",
  1107 => x"81c984c1",
  1108 => x"b7496997",
  1109 => x"87c204ac",
  1110 => x"976e4cc0",
  1111 => x"66c84abf",
  1112 => x"ff317249",
  1113 => x"9966c4b9",
  1114 => x"30724874",
  1115 => x"71484a70",
  1116 => x"ccdec2b0",
  1117 => x"d4e4c058",
  1118 => x"d449c087",
  1119 => x"497587c8",
  1120 => x"87c9f6c0",
  1121 => x"faf28ef4",
  1122 => x"1e731e87",
  1123 => x"fe494b71",
  1124 => x"497387cb",
  1125 => x"f287c6fe",
  1126 => x"731e87ed",
  1127 => x"c64b711e",
  1128 => x"db024aa3",
  1129 => x"028ac187",
  1130 => x"028a87d6",
  1131 => x"8a87dac1",
  1132 => x"87fcc002",
  1133 => x"e1c0028a",
  1134 => x"cb028a87",
  1135 => x"87dbc187",
  1136 => x"c7f649c7",
  1137 => x"87dec187",
  1138 => x"bfd8dac2",
  1139 => x"87cbc102",
  1140 => x"c288c148",
  1141 => x"c158dcda",
  1142 => x"dac287c1",
  1143 => x"c002bfdc",
  1144 => x"dac287f9",
  1145 => x"c148bfd8",
  1146 => x"dcdac280",
  1147 => x"87ebc058",
  1148 => x"bfd8dac2",
  1149 => x"c289c649",
  1150 => x"c059dcda",
  1151 => x"da03a9b7",
  1152 => x"d8dac287",
  1153 => x"d278c048",
  1154 => x"dcdac287",
  1155 => x"87cb02bf",
  1156 => x"bfd8dac2",
  1157 => x"c280c648",
  1158 => x"c058dcda",
  1159 => x"87e6d149",
  1160 => x"f3c04973",
  1161 => x"def087e7",
  1162 => x"5b5e0e87",
  1163 => x"ff0e5d5c",
  1164 => x"a6dc86d4",
  1165 => x"48a6c859",
  1166 => x"80c478c0",
  1167 => x"7866c0c1",
  1168 => x"78c180c4",
  1169 => x"78c180c4",
  1170 => x"48dcdac2",
  1171 => x"dac278c1",
  1172 => x"de48bfc0",
  1173 => x"87c905a8",
  1174 => x"cc87f8f4",
  1175 => x"e4cf58a6",
  1176 => x"87e3e487",
  1177 => x"e487c5e5",
  1178 => x"4c7087d2",
  1179 => x"02acfbc0",
  1180 => x"d887fbc1",
  1181 => x"edc10566",
  1182 => x"66fcc087",
  1183 => x"6a82c44a",
  1184 => x"c11e727e",
  1185 => x"c448fad9",
  1186 => x"a1c84966",
  1187 => x"7141204a",
  1188 => x"87f905aa",
  1189 => x"4a265110",
  1190 => x"4866fcc0",
  1191 => x"78dcc3c1",
  1192 => x"81c7496a",
  1193 => x"fcc05174",
  1194 => x"81c84966",
  1195 => x"fcc051c1",
  1196 => x"81c94966",
  1197 => x"fcc051c0",
  1198 => x"81ca4966",
  1199 => x"1ec151c0",
  1200 => x"496a1ed8",
  1201 => x"f7e381c8",
  1202 => x"c186c887",
  1203 => x"c04866c0",
  1204 => x"87c701a8",
  1205 => x"c148a6c8",
  1206 => x"c187ce78",
  1207 => x"c14866c0",
  1208 => x"58a6d088",
  1209 => x"c3e387c3",
  1210 => x"48a6d087",
  1211 => x"9c7478c2",
  1212 => x"87cdcd02",
  1213 => x"c14866c8",
  1214 => x"03a866c4",
  1215 => x"dc87c2cd",
  1216 => x"78c048a6",
  1217 => x"78c080e8",
  1218 => x"7087f1e1",
  1219 => x"acd0c14c",
  1220 => x"87d5c205",
  1221 => x"e47e66c4",
  1222 => x"a6c887d5",
  1223 => x"87dce158",
  1224 => x"ecc04c70",
  1225 => x"ebc105ac",
  1226 => x"4966c887",
  1227 => x"fcc091cb",
  1228 => x"a1c48166",
  1229 => x"c84d6a4a",
  1230 => x"66c44aa1",
  1231 => x"ccfdc052",
  1232 => x"87f8e079",
  1233 => x"029c4c70",
  1234 => x"fbc087d8",
  1235 => x"87d202ac",
  1236 => x"e7e05574",
  1237 => x"9c4c7087",
  1238 => x"c087c702",
  1239 => x"ff05acfb",
  1240 => x"e0c087ee",
  1241 => x"55c1c255",
  1242 => x"d87d97c0",
  1243 => x"a86e4866",
  1244 => x"c887db05",
  1245 => x"66cc4866",
  1246 => x"87ca04a8",
  1247 => x"c14866c8",
  1248 => x"58a6cc80",
  1249 => x"66cc87c8",
  1250 => x"d088c148",
  1251 => x"dfff58a6",
  1252 => x"4c7087ea",
  1253 => x"05acd0c1",
  1254 => x"66d487c8",
  1255 => x"d880c148",
  1256 => x"d0c158a6",
  1257 => x"ebfd02ac",
  1258 => x"4866c487",
  1259 => x"05a866d8",
  1260 => x"c087e0c9",
  1261 => x"c048a6e0",
  1262 => x"c0487478",
  1263 => x"7e7088fb",
  1264 => x"c9029848",
  1265 => x"cb4887e2",
  1266 => x"487e7088",
  1267 => x"cdc10298",
  1268 => x"88c94887",
  1269 => x"98487e70",
  1270 => x"87fec302",
  1271 => x"7088c448",
  1272 => x"0298487e",
  1273 => x"c14887ce",
  1274 => x"487e7088",
  1275 => x"e9c30298",
  1276 => x"87d6c887",
  1277 => x"c048a6dc",
  1278 => x"ddff78f0",
  1279 => x"4c7087fe",
  1280 => x"02acecc0",
  1281 => x"c087c4c0",
  1282 => x"c05ca6e0",
  1283 => x"cd02acec",
  1284 => x"e7ddff87",
  1285 => x"c04c7087",
  1286 => x"ff05acec",
  1287 => x"ecc087f3",
  1288 => x"c4c002ac",
  1289 => x"d3ddff87",
  1290 => x"ca1ec087",
  1291 => x"4966d01e",
  1292 => x"c4c191cb",
  1293 => x"80714866",
  1294 => x"c858a6cc",
  1295 => x"80c44866",
  1296 => x"cc58a6d0",
  1297 => x"ff49bf66",
  1298 => x"c187f5dd",
  1299 => x"d41ede1e",
  1300 => x"ff49bf66",
  1301 => x"d087e9dd",
  1302 => x"48497086",
  1303 => x"c08808c0",
  1304 => x"c058a6e8",
  1305 => x"eec006a8",
  1306 => x"66e4c087",
  1307 => x"03a8dd48",
  1308 => x"c487e4c0",
  1309 => x"c049bf66",
  1310 => x"c08166e4",
  1311 => x"e4c051e0",
  1312 => x"81c14966",
  1313 => x"81bf66c4",
  1314 => x"c051c1c2",
  1315 => x"c24966e4",
  1316 => x"bf66c481",
  1317 => x"6e51c081",
  1318 => x"dcc3c148",
  1319 => x"c8496e78",
  1320 => x"5166d081",
  1321 => x"81c9496e",
  1322 => x"6e5166d4",
  1323 => x"dc81ca49",
  1324 => x"66d05166",
  1325 => x"d480c148",
  1326 => x"66c858a6",
  1327 => x"a866cc48",
  1328 => x"87cbc004",
  1329 => x"c14866c8",
  1330 => x"58a6cc80",
  1331 => x"cc87d9c5",
  1332 => x"88c14866",
  1333 => x"c558a6d0",
  1334 => x"ddff87ce",
  1335 => x"e8c087d1",
  1336 => x"ddff58a6",
  1337 => x"e0c087c9",
  1338 => x"ecc058a6",
  1339 => x"cac005a8",
  1340 => x"48a6dc87",
  1341 => x"7866e4c0",
  1342 => x"ff87c4c0",
  1343 => x"c887fdd9",
  1344 => x"91cb4966",
  1345 => x"4866fcc0",
  1346 => x"7e708071",
  1347 => x"6e82c84a",
  1348 => x"c081ca49",
  1349 => x"dc5166e4",
  1350 => x"81c14966",
  1351 => x"8966e4c0",
  1352 => x"307148c1",
  1353 => x"89c14970",
  1354 => x"c27a9771",
  1355 => x"49bfc8de",
  1356 => x"2966e4c0",
  1357 => x"484a6a97",
  1358 => x"ecc09871",
  1359 => x"496e58a6",
  1360 => x"4d6981c4",
  1361 => x"c44866d8",
  1362 => x"c002a866",
  1363 => x"a6c487c8",
  1364 => x"c078c048",
  1365 => x"a6c487c5",
  1366 => x"c478c148",
  1367 => x"e0c01e66",
  1368 => x"ff49751e",
  1369 => x"c887d9d9",
  1370 => x"c04c7086",
  1371 => x"c106acb7",
  1372 => x"857487d4",
  1373 => x"7449e0c0",
  1374 => x"c14b7589",
  1375 => x"714ac3da",
  1376 => x"87e3ecfe",
  1377 => x"e0c085c2",
  1378 => x"80c14866",
  1379 => x"58a6e4c0",
  1380 => x"4966e8c0",
  1381 => x"a97081c1",
  1382 => x"87c8c002",
  1383 => x"c048a6c4",
  1384 => x"87c5c078",
  1385 => x"c148a6c4",
  1386 => x"1e66c478",
  1387 => x"c049a4c2",
  1388 => x"887148e0",
  1389 => x"751e4970",
  1390 => x"c3d8ff49",
  1391 => x"c086c887",
  1392 => x"ff01a8b7",
  1393 => x"e0c087c0",
  1394 => x"d1c00266",
  1395 => x"c9496e87",
  1396 => x"66e0c081",
  1397 => x"c1486e51",
  1398 => x"c078ddc4",
  1399 => x"496e87cc",
  1400 => x"51c281c9",
  1401 => x"c6c1486e",
  1402 => x"66c878c9",
  1403 => x"a866cc48",
  1404 => x"87cbc004",
  1405 => x"c14866c8",
  1406 => x"58a6cc80",
  1407 => x"cc87e9c0",
  1408 => x"88c14866",
  1409 => x"c058a6d0",
  1410 => x"d6ff87de",
  1411 => x"4c7087de",
  1412 => x"c187d5c0",
  1413 => x"c005acc6",
  1414 => x"66d087c8",
  1415 => x"d480c148",
  1416 => x"d6ff58a6",
  1417 => x"4c7087c6",
  1418 => x"c14866d4",
  1419 => x"58a6d880",
  1420 => x"c0029c74",
  1421 => x"66c887cb",
  1422 => x"66c4c148",
  1423 => x"fef204a8",
  1424 => x"ded5ff87",
  1425 => x"4866c887",
  1426 => x"c003a8c7",
  1427 => x"dac287e5",
  1428 => x"78c048dc",
  1429 => x"cb4966c8",
  1430 => x"66fcc091",
  1431 => x"4aa1c481",
  1432 => x"52c04a6a",
  1433 => x"4866c879",
  1434 => x"a6cc80c1",
  1435 => x"04a8c758",
  1436 => x"ff87dbff",
  1437 => x"dfff8ed4",
  1438 => x"6f4c87c9",
  1439 => x"2a206461",
  1440 => x"3a00202e",
  1441 => x"731e0020",
  1442 => x"9b4b711e",
  1443 => x"c287c602",
  1444 => x"c048d8da",
  1445 => x"c21ec778",
  1446 => x"1ebfd8da",
  1447 => x"1eefddc1",
  1448 => x"bfc0dac2",
  1449 => x"87c1ee49",
  1450 => x"dac286cc",
  1451 => x"e249bfc0",
  1452 => x"9b7387f9",
  1453 => x"c187c802",
  1454 => x"c049efdd",
  1455 => x"ff87e0e2",
  1456 => x"1e87c4de",
  1457 => x"48dbddc1",
  1458 => x"dfc150c0",
  1459 => x"ff49bfd2",
  1460 => x"c087e4d8",
  1461 => x"1e4f2648",
  1462 => x"c187dbc7",
  1463 => x"87e6fe49",
  1464 => x"87cceffe",
  1465 => x"cd029870",
  1466 => x"e6f6fe87",
  1467 => x"02987087",
  1468 => x"4ac187c4",
  1469 => x"4ac087c2",
  1470 => x"ce059a72",
  1471 => x"c11ec087",
  1472 => x"c049f2dc",
  1473 => x"c487dbee",
  1474 => x"c287fe86",
  1475 => x"c048d8da",
  1476 => x"c0dac278",
  1477 => x"1e78c048",
  1478 => x"49fddcc1",
  1479 => x"87c2eec0",
  1480 => x"defe1ec0",
  1481 => x"c0497087",
  1482 => x"c387f7ed",
  1483 => x"8ef887c7",
  1484 => x"44534f26",
  1485 => x"69616620",
  1486 => x"2e64656c",
  1487 => x"6f6f4200",
  1488 => x"676e6974",
  1489 => x"002e2e2e",
  1490 => x"cfe2c01e",
  1491 => x"2687fa87",
  1492 => x"c2fe1e4f",
  1493 => x"c087f187",
  1494 => x"004f2648",
  1495 => x"00000100",
  1496 => x"45208000",
  1497 => x"00746978",
  1498 => x"61422080",
  1499 => x"99006b63",
  1500 => x"ac00000e",
  1501 => x"00000026",
  1502 => x"0e990000",
  1503 => x"26ca0000",
  1504 => x"00000000",
  1505 => x"000e9900",
  1506 => x"0026e800",
  1507 => x"00000000",
  1508 => x"00000e99",
  1509 => x"00002706",
  1510 => x"99000000",
  1511 => x"2400000e",
  1512 => x"00000027",
  1513 => x"0e990000",
  1514 => x"27420000",
  1515 => x"00000000",
  1516 => x"000e9900",
  1517 => x"00276000",
  1518 => x"00000000",
  1519 => x"00000f4c",
  1520 => x"00000000",
  1521 => x"9a000000",
  1522 => x"00000011",
  1523 => x"00000000",
  1524 => x"17d60000",
  1525 => x"4f420000",
  1526 => x"2020544f",
  1527 => x"4f522020",
  1528 => x"fe1e004d",
  1529 => x"78c048f0",
  1530 => x"097909cd",
  1531 => x"fe1e4f26",
  1532 => x"2648bff0",
  1533 => x"f0fe1e4f",
  1534 => x"2678c148",
  1535 => x"f0fe1e4f",
  1536 => x"2678c048",
  1537 => x"4a711e4f",
  1538 => x"265252c0",
  1539 => x"5b5e0e4f",
  1540 => x"f40e5d5c",
  1541 => x"974d7186",
  1542 => x"a5c17e6d",
  1543 => x"486c974c",
  1544 => x"6e58a6c8",
  1545 => x"a866c448",
  1546 => x"ff87c505",
  1547 => x"87e6c048",
  1548 => x"c287caff",
  1549 => x"6c9749a5",
  1550 => x"4ba3714b",
  1551 => x"974b6b97",
  1552 => x"486e7e6c",
  1553 => x"a6c880c1",
  1554 => x"cc98c758",
  1555 => x"977058a6",
  1556 => x"87e1fe7c",
  1557 => x"8ef44873",
  1558 => x"4c264d26",
  1559 => x"4f264b26",
  1560 => x"5c5b5e0e",
  1561 => x"7186f40e",
  1562 => x"4a66d84c",
  1563 => x"c29affc3",
  1564 => x"6c974ba4",
  1565 => x"49a17349",
  1566 => x"6c975172",
  1567 => x"c1486e7e",
  1568 => x"58a6c880",
  1569 => x"a6cc98c7",
  1570 => x"f4547058",
  1571 => x"87caff8e",
  1572 => x"e8fd1e1e",
  1573 => x"4abfe087",
  1574 => x"c0e0c049",
  1575 => x"87cb0299",
  1576 => x"ddc21e72",
  1577 => x"f7fe49fe",
  1578 => x"fd86c487",
  1579 => x"7e7087c0",
  1580 => x"2687c2fd",
  1581 => x"c21e4f26",
  1582 => x"fd49fedd",
  1583 => x"e2c187c7",
  1584 => x"ddfc49d0",
  1585 => x"87eec387",
  1586 => x"5e0e4f26",
  1587 => x"0e5d5c5b",
  1588 => x"ddc24d71",
  1589 => x"f4fc49fe",
  1590 => x"c04b7087",
  1591 => x"c304abb7",
  1592 => x"f0c387c2",
  1593 => x"87c905ab",
  1594 => x"48eee6c1",
  1595 => x"e3c278c1",
  1596 => x"abe0c387",
  1597 => x"c187c905",
  1598 => x"c148f2e6",
  1599 => x"87d4c278",
  1600 => x"bff2e6c1",
  1601 => x"c287c602",
  1602 => x"c24ca3c0",
  1603 => x"c14c7387",
  1604 => x"02bfeee6",
  1605 => x"7487e0c0",
  1606 => x"29b7c449",
  1607 => x"c5e8c191",
  1608 => x"cf4a7481",
  1609 => x"c192c29a",
  1610 => x"70307248",
  1611 => x"72baff4a",
  1612 => x"70986948",
  1613 => x"7487db79",
  1614 => x"29b7c449",
  1615 => x"c5e8c191",
  1616 => x"cf4a7481",
  1617 => x"c392c29a",
  1618 => x"70307248",
  1619 => x"b069484a",
  1620 => x"9d757970",
  1621 => x"87f0c005",
  1622 => x"c848d0ff",
  1623 => x"d4ff78e1",
  1624 => x"c178c548",
  1625 => x"02bff2e6",
  1626 => x"e0c387c3",
  1627 => x"eee6c178",
  1628 => x"87c602bf",
  1629 => x"c348d4ff",
  1630 => x"d4ff78f0",
  1631 => x"ff0b7b0b",
  1632 => x"e1c848d0",
  1633 => x"78e0c078",
  1634 => x"48f2e6c1",
  1635 => x"e6c178c0",
  1636 => x"78c048ee",
  1637 => x"49feddc2",
  1638 => x"7087f2f9",
  1639 => x"abb7c04b",
  1640 => x"87fefc03",
  1641 => x"4d2648c0",
  1642 => x"4b264c26",
  1643 => x"00004f26",
  1644 => x"00000000",
  1645 => x"c01e0000",
  1646 => x"c449724a",
  1647 => x"c5e8c191",
  1648 => x"c179c081",
  1649 => x"aab7d082",
  1650 => x"2687ee04",
  1651 => x"5b5e0e4f",
  1652 => x"710e5d5c",
  1653 => x"87e5f84d",
  1654 => x"b7c44a75",
  1655 => x"e8c1922a",
  1656 => x"4c7582c5",
  1657 => x"94c29ccf",
  1658 => x"744b496a",
  1659 => x"c29bc32b",
  1660 => x"70307448",
  1661 => x"74bcff4c",
  1662 => x"70987148",
  1663 => x"87f5f77a",
  1664 => x"e1fe4873",
  1665 => x"00000087",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"d0ff1e00",
  1682 => x"78e1c848",
  1683 => x"d4ff4871",
  1684 => x"66c47808",
  1685 => x"08d4ff48",
  1686 => x"1e4f2678",
  1687 => x"66c44a71",
  1688 => x"49721e49",
  1689 => x"ff87deff",
  1690 => x"e0c048d0",
  1691 => x"4f262678",
  1692 => x"711e731e",
  1693 => x"4966c84b",
  1694 => x"c14a731e",
  1695 => x"ff49a2e0",
  1696 => x"c42687d9",
  1697 => x"264d2687",
  1698 => x"264b264c",
  1699 => x"d4ff1e4f",
  1700 => x"7affc34a",
  1701 => x"c048d0ff",
  1702 => x"7ade78e1",
  1703 => x"bfc8dec2",
  1704 => x"c848497a",
  1705 => x"717a7028",
  1706 => x"7028d048",
  1707 => x"d848717a",
  1708 => x"ff7a7028",
  1709 => x"e0c048d0",
  1710 => x"1e4f2678",
  1711 => x"c848d0ff",
  1712 => x"487178c9",
  1713 => x"7808d4ff",
  1714 => x"711e4f26",
  1715 => x"87eb494a",
  1716 => x"c848d0ff",
  1717 => x"1e4f2678",
  1718 => x"4b711e73",
  1719 => x"bfd8dec2",
  1720 => x"c287c302",
  1721 => x"d0ff87eb",
  1722 => x"78c9c848",
  1723 => x"e0c04873",
  1724 => x"08d4ffb0",
  1725 => x"ccdec278",
  1726 => x"c878c048",
  1727 => x"87c50266",
  1728 => x"c249ffc3",
  1729 => x"c249c087",
  1730 => x"cc59d4de",
  1731 => x"87c60266",
  1732 => x"4ad5d5c5",
  1733 => x"ffcf87c4",
  1734 => x"dec24aff",
  1735 => x"dec25ad8",
  1736 => x"78c148d8",
  1737 => x"4d2687c4",
  1738 => x"4b264c26",
  1739 => x"5e0e4f26",
  1740 => x"0e5d5c5b",
  1741 => x"dec24a71",
  1742 => x"724cbfd4",
  1743 => x"87cb029a",
  1744 => x"c191c849",
  1745 => x"714bcdeb",
  1746 => x"c187c483",
  1747 => x"c04bcdef",
  1748 => x"7449134d",
  1749 => x"d0dec299",
  1750 => x"b87148bf",
  1751 => x"7808d4ff",
  1752 => x"852cb7c1",
  1753 => x"04adb7c8",
  1754 => x"dec287e7",
  1755 => x"c848bfcc",
  1756 => x"d0dec280",
  1757 => x"87eefe58",
  1758 => x"711e731e",
  1759 => x"9a4a134b",
  1760 => x"7287cb02",
  1761 => x"87e6fe49",
  1762 => x"059a4a13",
  1763 => x"d9fe87f5",
  1764 => x"dec21e87",
  1765 => x"c249bfcc",
  1766 => x"c148ccde",
  1767 => x"c0c478a1",
  1768 => x"db03a9b7",
  1769 => x"48d4ff87",
  1770 => x"bfd0dec2",
  1771 => x"ccdec278",
  1772 => x"dec249bf",
  1773 => x"a1c148cc",
  1774 => x"b7c0c478",
  1775 => x"87e504a9",
  1776 => x"c848d0ff",
  1777 => x"d8dec278",
  1778 => x"2678c048",
  1779 => x"0000004f",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00005f5f",
  1783 => x"03030000",
  1784 => x"00030300",
  1785 => x"7f7f1400",
  1786 => x"147f7f14",
  1787 => x"2e240000",
  1788 => x"123a6b6b",
  1789 => x"366a4c00",
  1790 => x"32566c18",
  1791 => x"4f7e3000",
  1792 => x"683a7759",
  1793 => x"04000040",
  1794 => x"00000307",
  1795 => x"1c000000",
  1796 => x"0041633e",
  1797 => x"41000000",
  1798 => x"001c3e63",
  1799 => x"3e2a0800",
  1800 => x"2a3e1c1c",
  1801 => x"08080008",
  1802 => x"08083e3e",
  1803 => x"80000000",
  1804 => x"000060e0",
  1805 => x"08080000",
  1806 => x"08080808",
  1807 => x"00000000",
  1808 => x"00006060",
  1809 => x"30604000",
  1810 => x"03060c18",
  1811 => x"7f3e0001",
  1812 => x"3e7f4d59",
  1813 => x"06040000",
  1814 => x"00007f7f",
  1815 => x"63420000",
  1816 => x"464f5971",
  1817 => x"63220000",
  1818 => x"367f4949",
  1819 => x"161c1800",
  1820 => x"107f7f13",
  1821 => x"67270000",
  1822 => x"397d4545",
  1823 => x"7e3c0000",
  1824 => x"3079494b",
  1825 => x"01010000",
  1826 => x"070f7971",
  1827 => x"7f360000",
  1828 => x"367f4949",
  1829 => x"4f060000",
  1830 => x"1e3f6949",
  1831 => x"00000000",
  1832 => x"00006666",
  1833 => x"80000000",
  1834 => x"000066e6",
  1835 => x"08080000",
  1836 => x"22221414",
  1837 => x"14140000",
  1838 => x"14141414",
  1839 => x"22220000",
  1840 => x"08081414",
  1841 => x"03020000",
  1842 => x"060f5951",
  1843 => x"417f3e00",
  1844 => x"1e1f555d",
  1845 => x"7f7e0000",
  1846 => x"7e7f0909",
  1847 => x"7f7f0000",
  1848 => x"367f4949",
  1849 => x"3e1c0000",
  1850 => x"41414163",
  1851 => x"7f7f0000",
  1852 => x"1c3e6341",
  1853 => x"7f7f0000",
  1854 => x"41414949",
  1855 => x"7f7f0000",
  1856 => x"01010909",
  1857 => x"7f3e0000",
  1858 => x"7a7b4941",
  1859 => x"7f7f0000",
  1860 => x"7f7f0808",
  1861 => x"41000000",
  1862 => x"00417f7f",
  1863 => x"60200000",
  1864 => x"3f7f4040",
  1865 => x"087f7f00",
  1866 => x"4163361c",
  1867 => x"7f7f0000",
  1868 => x"40404040",
  1869 => x"067f7f00",
  1870 => x"7f7f060c",
  1871 => x"067f7f00",
  1872 => x"7f7f180c",
  1873 => x"7f3e0000",
  1874 => x"3e7f4141",
  1875 => x"7f7f0000",
  1876 => x"060f0909",
  1877 => x"417f3e00",
  1878 => x"407e7f61",
  1879 => x"7f7f0000",
  1880 => x"667f1909",
  1881 => x"6f260000",
  1882 => x"327b594d",
  1883 => x"01010000",
  1884 => x"01017f7f",
  1885 => x"7f3f0000",
  1886 => x"3f7f4040",
  1887 => x"3f0f0000",
  1888 => x"0f3f7070",
  1889 => x"307f7f00",
  1890 => x"7f7f3018",
  1891 => x"36634100",
  1892 => x"63361c1c",
  1893 => x"06030141",
  1894 => x"03067c7c",
  1895 => x"59716101",
  1896 => x"4143474d",
  1897 => x"7f000000",
  1898 => x"0041417f",
  1899 => x"06030100",
  1900 => x"6030180c",
  1901 => x"41000040",
  1902 => x"007f7f41",
  1903 => x"060c0800",
  1904 => x"080c0603",
  1905 => x"80808000",
  1906 => x"80808080",
  1907 => x"00000000",
  1908 => x"00040703",
  1909 => x"74200000",
  1910 => x"787c5454",
  1911 => x"7f7f0000",
  1912 => x"387c4444",
  1913 => x"7c380000",
  1914 => x"00444444",
  1915 => x"7c380000",
  1916 => x"7f7f4444",
  1917 => x"7c380000",
  1918 => x"185c5454",
  1919 => x"7e040000",
  1920 => x"0005057f",
  1921 => x"bc180000",
  1922 => x"7cfca4a4",
  1923 => x"7f7f0000",
  1924 => x"787c0404",
  1925 => x"00000000",
  1926 => x"00407d3d",
  1927 => x"80800000",
  1928 => x"007dfd80",
  1929 => x"7f7f0000",
  1930 => x"446c3810",
  1931 => x"00000000",
  1932 => x"00407f3f",
  1933 => x"0c7c7c00",
  1934 => x"787c0c18",
  1935 => x"7c7c0000",
  1936 => x"787c0404",
  1937 => x"7c380000",
  1938 => x"387c4444",
  1939 => x"fcfc0000",
  1940 => x"183c2424",
  1941 => x"3c180000",
  1942 => x"fcfc2424",
  1943 => x"7c7c0000",
  1944 => x"080c0404",
  1945 => x"5c480000",
  1946 => x"20745454",
  1947 => x"3f040000",
  1948 => x"0044447f",
  1949 => x"7c3c0000",
  1950 => x"7c7c4040",
  1951 => x"3c1c0000",
  1952 => x"1c3c6060",
  1953 => x"607c3c00",
  1954 => x"3c7c6030",
  1955 => x"386c4400",
  1956 => x"446c3810",
  1957 => x"bc1c0000",
  1958 => x"1c3c60e0",
  1959 => x"64440000",
  1960 => x"444c5c74",
  1961 => x"08080000",
  1962 => x"4141773e",
  1963 => x"00000000",
  1964 => x"00007f7f",
  1965 => x"41410000",
  1966 => x"08083e77",
  1967 => x"01010200",
  1968 => x"01020203",
  1969 => x"7f7f7f00",
  1970 => x"7f7f7f7f",
  1971 => x"1c080800",
  1972 => x"7f3e3e1c",
  1973 => x"3e7f7f7f",
  1974 => x"081c1c3e",
  1975 => x"18100008",
  1976 => x"10187c7c",
  1977 => x"30100000",
  1978 => x"10307c7c",
  1979 => x"60301000",
  1980 => x"061e7860",
  1981 => x"3c664200",
  1982 => x"42663c18",
  1983 => x"6a387800",
  1984 => x"386cc6c2",
  1985 => x"00006000",
  1986 => x"60000060",
  1987 => x"5b5e0e00",
  1988 => x"1e0e5d5c",
  1989 => x"dec24c71",
  1990 => x"c04dbfdd",
  1991 => x"741ec04b",
  1992 => x"87c702ab",
  1993 => x"c048a6c4",
  1994 => x"c487c578",
  1995 => x"78c148a6",
  1996 => x"731e66c4",
  1997 => x"87dfee49",
  1998 => x"e0c086c8",
  1999 => x"87eeef49",
  2000 => x"6a4aa5c4",
  2001 => x"87f0f049",
  2002 => x"cb87c6f1",
  2003 => x"c883c185",
  2004 => x"ff04abb7",
  2005 => x"262687c7",
  2006 => x"264c264d",
  2007 => x"1e4f264b",
  2008 => x"dec24a71",
  2009 => x"dec25ae1",
  2010 => x"78c748e1",
  2011 => x"87ddfe49",
  2012 => x"731e4f26",
  2013 => x"c04a711e",
  2014 => x"d303aab7",
  2015 => x"fbcbc287",
  2016 => x"87c405bf",
  2017 => x"87c24bc1",
  2018 => x"cbc24bc0",
  2019 => x"87c45bff",
  2020 => x"5affcbc2",
  2021 => x"bffbcbc2",
  2022 => x"c19ac14a",
  2023 => x"ec49a2c0",
  2024 => x"48fc87e8",
  2025 => x"bffbcbc2",
  2026 => x"87effe78",
  2027 => x"c44a711e",
  2028 => x"49721e66",
  2029 => x"2687f9ea",
  2030 => x"ff1e4f26",
  2031 => x"ffc348d4",
  2032 => x"48d0ff78",
  2033 => x"ff78e1c0",
  2034 => x"78c148d4",
  2035 => x"30c44871",
  2036 => x"7808d4ff",
  2037 => x"c048d0ff",
  2038 => x"4f2678e0",
  2039 => x"5c5b5e0e",
  2040 => x"86f00e5d",
  2041 => x"c048a6c8",
  2042 => x"ec4b4d78",
  2043 => x"80fc7ebf",
  2044 => x"bfdddec2",
  2045 => x"4cbfe878",
  2046 => x"bffbcbc2",
  2047 => x"87cae349",
  2048 => x"cb49eecb",
  2049 => x"a6d087fd",
  2050 => x"e649c758",
  2051 => x"987087ff",
  2052 => x"6e87c805",
  2053 => x"0299c149",
  2054 => x"c187c3c1",
  2055 => x"7ebfec4b",
  2056 => x"bffbcbc2",
  2057 => x"87e2e249",
  2058 => x"cb4966cc",
  2059 => x"987087e1",
  2060 => x"c287d802",
  2061 => x"49bff3cb",
  2062 => x"cbc2b9c1",
  2063 => x"fd7159f7",
  2064 => x"eecb87f8",
  2065 => x"87fbca49",
  2066 => x"c758a6d0",
  2067 => x"87fde549",
  2068 => x"ff059870",
  2069 => x"496e87c5",
  2070 => x"fe0599c1",
  2071 => x"9b7387fd",
  2072 => x"ff87d002",
  2073 => x"87cafc49",
  2074 => x"e549dac1",
  2075 => x"a6c887df",
  2076 => x"c278c148",
  2077 => x"05bffbcb",
  2078 => x"c387e9c0",
  2079 => x"cce549fd",
  2080 => x"49fac387",
  2081 => x"7487c6e5",
  2082 => x"99ffc349",
  2083 => x"49c01e71",
  2084 => x"7487d9fc",
  2085 => x"29b7c849",
  2086 => x"49c11e71",
  2087 => x"c887cdfc",
  2088 => x"87f9c786",
  2089 => x"ffc34974",
  2090 => x"2cb7c899",
  2091 => x"9c74b471",
  2092 => x"c287dd02",
  2093 => x"49bff7cb",
  2094 => x"7087d4c9",
  2095 => x"87c40598",
  2096 => x"87d24cc0",
  2097 => x"c849e0c2",
  2098 => x"cbc287f9",
  2099 => x"87c658fb",
  2100 => x"48f7cbc2",
  2101 => x"497478c0",
  2102 => x"ce0599c2",
  2103 => x"49ebc387",
  2104 => x"7087eae3",
  2105 => x"0299c249",
  2106 => x"fb87c2c0",
  2107 => x"c149744d",
  2108 => x"87ce0599",
  2109 => x"e349f4c3",
  2110 => x"497087d3",
  2111 => x"c00299c2",
  2112 => x"4dfa87c2",
  2113 => x"99c84974",
  2114 => x"c387cd05",
  2115 => x"fce249f5",
  2116 => x"c2497087",
  2117 => x"87d90299",
  2118 => x"bfe1dec2",
  2119 => x"87cac002",
  2120 => x"c288c148",
  2121 => x"c058e5de",
  2122 => x"4dff87c2",
  2123 => x"c148a6c8",
  2124 => x"c4497478",
  2125 => x"cdc00599",
  2126 => x"49f2c387",
  2127 => x"7087cee2",
  2128 => x"0299c249",
  2129 => x"dec287df",
  2130 => x"487ebfe1",
  2131 => x"03a8b7c7",
  2132 => x"6e87cbc0",
  2133 => x"c280c148",
  2134 => x"c058e5de",
  2135 => x"4dfe87c2",
  2136 => x"c148a6c8",
  2137 => x"49fdc378",
  2138 => x"7087e2e1",
  2139 => x"0299c249",
  2140 => x"c287d8c0",
  2141 => x"02bfe1de",
  2142 => x"c287c9c0",
  2143 => x"c048e1de",
  2144 => x"87c2c078",
  2145 => x"a6c84dfd",
  2146 => x"c378c148",
  2147 => x"fce049fa",
  2148 => x"c2497087",
  2149 => x"dcc00299",
  2150 => x"e1dec287",
  2151 => x"b7c748bf",
  2152 => x"c9c003a8",
  2153 => x"e1dec287",
  2154 => x"c078c748",
  2155 => x"4dfc87c2",
  2156 => x"c148a6c8",
  2157 => x"adb7c078",
  2158 => x"87d0c003",
  2159 => x"c14a66c4",
  2160 => x"026a82d8",
  2161 => x"4b87c5c0",
  2162 => x"0f734975",
  2163 => x"dec24bc0",
  2164 => x"50c048dc",
  2165 => x"c449eecb",
  2166 => x"a6d087e9",
  2167 => x"dcdec258",
  2168 => x"c105bf97",
  2169 => x"497487de",
  2170 => x"0599f0c3",
  2171 => x"c187cdc0",
  2172 => x"dfff49da",
  2173 => x"987087d7",
  2174 => x"87c8c102",
  2175 => x"bfe84bc1",
  2176 => x"ffc3494c",
  2177 => x"2cb7c899",
  2178 => x"cbc2b471",
  2179 => x"ff49bffb",
  2180 => x"cc87f7da",
  2181 => x"f6c34966",
  2182 => x"02987087",
  2183 => x"c287c6c0",
  2184 => x"c148dcde",
  2185 => x"dcdec250",
  2186 => x"c005bf97",
  2187 => x"497487d6",
  2188 => x"0599f0c3",
  2189 => x"c187c5ff",
  2190 => x"deff49da",
  2191 => x"987087cf",
  2192 => x"87f8fe05",
  2193 => x"c0029b73",
  2194 => x"a6cc87e0",
  2195 => x"e1dec248",
  2196 => x"66cc78bf",
  2197 => x"c491cb49",
  2198 => x"80714866",
  2199 => x"bf6e7e70",
  2200 => x"87c6c002",
  2201 => x"4966cc4b",
  2202 => x"66c80f73",
  2203 => x"87c8c002",
  2204 => x"bfe1dec2",
  2205 => x"87d5f249",
  2206 => x"bfffcbc2",
  2207 => x"87ddc002",
  2208 => x"87cbc249",
  2209 => x"c0029870",
  2210 => x"dec287d3",
  2211 => x"f149bfe1",
  2212 => x"49c087fb",
  2213 => x"c287dbf3",
  2214 => x"c048ffcb",
  2215 => x"f28ef078",
  2216 => x"5e0e87f5",
  2217 => x"0e5d5c5b",
  2218 => x"c24c711e",
  2219 => x"49bfddde",
  2220 => x"4da1cdc1",
  2221 => x"6981d1c1",
  2222 => x"029c747e",
  2223 => x"a5c487cf",
  2224 => x"c27b744b",
  2225 => x"49bfddde",
  2226 => x"6e87d4f2",
  2227 => x"059c747b",
  2228 => x"4bc087c4",
  2229 => x"4bc187c2",
  2230 => x"d5f24973",
  2231 => x"0266d487",
  2232 => x"de4987c7",
  2233 => x"c24a7087",
  2234 => x"c24ac087",
  2235 => x"265ac3cc",
  2236 => x"0087e4f1",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"1e000000",
  2241 => x"c8ff4a71",
  2242 => x"a17249bf",
  2243 => x"1e4f2648",
  2244 => x"89bfc8ff",
  2245 => x"c0c0c0fe",
  2246 => x"01a9c0c0",
  2247 => x"4ac087c4",
  2248 => x"4ac187c2",
  2249 => x"4f264872",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
