
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"de",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f0",x"de",x"c2"),
    14 => (x"48",x"f0",x"cc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"cb",x"dc"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"48",x"72",x"4c"),
    72 => (x"7c",x"70",x"98",x"ff"),
    73 => (x"bf",x"f0",x"cc",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"ff",x"c3",x"48",x"71"),
    79 => (x"d0",x"7c",x"70",x"98"),
    80 => (x"29",x"d0",x"49",x"66"),
    81 => (x"ff",x"c3",x"48",x"71"),
    82 => (x"d0",x"7c",x"70",x"98"),
    83 => (x"29",x"c8",x"49",x"66"),
    84 => (x"ff",x"c3",x"48",x"71"),
    85 => (x"d0",x"7c",x"70",x"98"),
    86 => (x"ff",x"c3",x"48",x"66"),
    87 => (x"72",x"7c",x"70",x"98"),
    88 => (x"71",x"29",x"d0",x"49"),
    89 => (x"98",x"ff",x"c3",x"48"),
    90 => (x"4b",x"6c",x"7c",x"70"),
    91 => (x"4d",x"ff",x"f0",x"c9"),
    92 => (x"05",x"ab",x"ff",x"c3"),
    93 => (x"ff",x"c3",x"87",x"d0"),
    94 => (x"c1",x"4b",x"6c",x"7c"),
    95 => (x"87",x"c6",x"02",x"8d"),
    96 => (x"02",x"ab",x"ff",x"c3"),
    97 => (x"48",x"73",x"87",x"f0"),
    98 => (x"1e",x"87",x"ff",x"fd"),
    99 => (x"d4",x"ff",x"49",x"c0"),
   100 => (x"78",x"ff",x"c3",x"48"),
   101 => (x"c8",x"c3",x"81",x"c1"),
   102 => (x"f1",x"04",x"a9",x"b7"),
   103 => (x"1e",x"4f",x"26",x"87"),
   104 => (x"87",x"e7",x"1e",x"73"),
   105 => (x"4b",x"df",x"f8",x"c4"),
   106 => (x"ff",x"c0",x"1e",x"c0"),
   107 => (x"49",x"f7",x"c1",x"f0"),
   108 => (x"c4",x"87",x"df",x"fd"),
   109 => (x"05",x"a8",x"c1",x"86"),
   110 => (x"ff",x"87",x"ea",x"c0"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c0",x"c0",x"c1",x"78"),
   113 => (x"1e",x"c0",x"c0",x"c0"),
   114 => (x"c1",x"f0",x"e1",x"c0"),
   115 => (x"c1",x"fd",x"49",x"e9"),
   116 => (x"70",x"86",x"c4",x"87"),
   117 => (x"87",x"ca",x"05",x"98"),
   118 => (x"c3",x"48",x"d4",x"ff"),
   119 => (x"48",x"c1",x"78",x"ff"),
   120 => (x"e6",x"fe",x"87",x"cb"),
   121 => (x"05",x"8b",x"c1",x"87"),
   122 => (x"c0",x"87",x"fd",x"fe"),
   123 => (x"87",x"de",x"fc",x"48"),
   124 => (x"ff",x"1e",x"73",x"1e"),
   125 => (x"ff",x"c3",x"48",x"d4"),
   126 => (x"c0",x"4b",x"d3",x"78"),
   127 => (x"f0",x"ff",x"c0",x"1e"),
   128 => (x"fc",x"49",x"c1",x"c1"),
   129 => (x"86",x"c4",x"87",x"cc"),
   130 => (x"ca",x"05",x"98",x"70"),
   131 => (x"48",x"d4",x"ff",x"87"),
   132 => (x"c1",x"78",x"ff",x"c3"),
   133 => (x"fd",x"87",x"cb",x"48"),
   134 => (x"8b",x"c1",x"87",x"f1"),
   135 => (x"87",x"db",x"ff",x"05"),
   136 => (x"e9",x"fb",x"48",x"c0"),
   137 => (x"5b",x"5e",x"0e",x"87"),
   138 => (x"d4",x"ff",x"0e",x"5c"),
   139 => (x"87",x"db",x"fd",x"4c"),
   140 => (x"c0",x"1e",x"ea",x"c6"),
   141 => (x"c8",x"c1",x"f0",x"e1"),
   142 => (x"87",x"d6",x"fb",x"49"),
   143 => (x"a8",x"c1",x"86",x"c4"),
   144 => (x"fe",x"87",x"c8",x"02"),
   145 => (x"48",x"c0",x"87",x"ea"),
   146 => (x"fa",x"87",x"e2",x"c1"),
   147 => (x"49",x"70",x"87",x"d2"),
   148 => (x"99",x"ff",x"ff",x"cf"),
   149 => (x"02",x"a9",x"ea",x"c6"),
   150 => (x"d3",x"fe",x"87",x"c8"),
   151 => (x"c1",x"48",x"c0",x"87"),
   152 => (x"ff",x"c3",x"87",x"cb"),
   153 => (x"4b",x"f1",x"c0",x"7c"),
   154 => (x"70",x"87",x"f4",x"fc"),
   155 => (x"eb",x"c0",x"02",x"98"),
   156 => (x"c0",x"1e",x"c0",x"87"),
   157 => (x"fa",x"c1",x"f0",x"ff"),
   158 => (x"87",x"d6",x"fa",x"49"),
   159 => (x"98",x"70",x"86",x"c4"),
   160 => (x"c3",x"87",x"d9",x"05"),
   161 => (x"49",x"6c",x"7c",x"ff"),
   162 => (x"7c",x"7c",x"ff",x"c3"),
   163 => (x"c0",x"c1",x"7c",x"7c"),
   164 => (x"87",x"c4",x"02",x"99"),
   165 => (x"87",x"d5",x"48",x"c1"),
   166 => (x"87",x"d1",x"48",x"c0"),
   167 => (x"c4",x"05",x"ab",x"c2"),
   168 => (x"c8",x"48",x"c0",x"87"),
   169 => (x"05",x"8b",x"c1",x"87"),
   170 => (x"c0",x"87",x"fd",x"fe"),
   171 => (x"87",x"dc",x"f9",x"48"),
   172 => (x"c2",x"1e",x"73",x"1e"),
   173 => (x"c1",x"48",x"f0",x"cc"),
   174 => (x"ff",x"4b",x"c7",x"78"),
   175 => (x"78",x"c2",x"48",x"d0"),
   176 => (x"ff",x"87",x"c8",x"fb"),
   177 => (x"78",x"c3",x"48",x"d0"),
   178 => (x"e5",x"c0",x"1e",x"c0"),
   179 => (x"49",x"c0",x"c1",x"d0"),
   180 => (x"c4",x"87",x"ff",x"f8"),
   181 => (x"05",x"a8",x"c1",x"86"),
   182 => (x"c2",x"4b",x"87",x"c1"),
   183 => (x"87",x"c5",x"05",x"ab"),
   184 => (x"f9",x"c0",x"48",x"c0"),
   185 => (x"05",x"8b",x"c1",x"87"),
   186 => (x"fc",x"87",x"d0",x"ff"),
   187 => (x"cc",x"c2",x"87",x"f7"),
   188 => (x"98",x"70",x"58",x"f4"),
   189 => (x"c1",x"87",x"cd",x"05"),
   190 => (x"f0",x"ff",x"c0",x"1e"),
   191 => (x"f8",x"49",x"d0",x"c1"),
   192 => (x"86",x"c4",x"87",x"d0"),
   193 => (x"c3",x"48",x"d4",x"ff"),
   194 => (x"fd",x"c2",x"78",x"ff"),
   195 => (x"f8",x"cc",x"c2",x"87"),
   196 => (x"48",x"d0",x"ff",x"58"),
   197 => (x"d4",x"ff",x"78",x"c2"),
   198 => (x"78",x"ff",x"c3",x"48"),
   199 => (x"ed",x"f7",x"48",x"c1"),
   200 => (x"5b",x"5e",x"0e",x"87"),
   201 => (x"71",x"0e",x"5d",x"5c"),
   202 => (x"c5",x"4c",x"c0",x"4b"),
   203 => (x"4a",x"df",x"cd",x"ee"),
   204 => (x"c3",x"48",x"d4",x"ff"),
   205 => (x"48",x"68",x"78",x"ff"),
   206 => (x"05",x"a8",x"fe",x"c3"),
   207 => (x"ff",x"87",x"fe",x"c0"),
   208 => (x"9b",x"73",x"4d",x"d4"),
   209 => (x"d0",x"87",x"cc",x"02"),
   210 => (x"49",x"73",x"1e",x"66"),
   211 => (x"c4",x"87",x"e8",x"f5"),
   212 => (x"ff",x"87",x"d6",x"86"),
   213 => (x"d1",x"c4",x"48",x"d0"),
   214 => (x"7d",x"ff",x"c3",x"78"),
   215 => (x"c1",x"48",x"66",x"d0"),
   216 => (x"58",x"a6",x"d4",x"88"),
   217 => (x"f0",x"05",x"98",x"70"),
   218 => (x"48",x"d4",x"ff",x"87"),
   219 => (x"78",x"78",x"ff",x"c3"),
   220 => (x"c5",x"05",x"9b",x"73"),
   221 => (x"48",x"d0",x"ff",x"87"),
   222 => (x"4a",x"c1",x"78",x"d0"),
   223 => (x"05",x"8a",x"c1",x"4c"),
   224 => (x"74",x"87",x"ed",x"fe"),
   225 => (x"87",x"c2",x"f6",x"48"),
   226 => (x"71",x"1e",x"73",x"1e"),
   227 => (x"ff",x"4b",x"c0",x"4a"),
   228 => (x"ff",x"c3",x"48",x"d4"),
   229 => (x"48",x"d0",x"ff",x"78"),
   230 => (x"ff",x"78",x"c3",x"c4"),
   231 => (x"ff",x"c3",x"48",x"d4"),
   232 => (x"c0",x"1e",x"72",x"78"),
   233 => (x"d1",x"c1",x"f0",x"ff"),
   234 => (x"87",x"e6",x"f5",x"49"),
   235 => (x"98",x"70",x"86",x"c4"),
   236 => (x"c8",x"87",x"d2",x"05"),
   237 => (x"66",x"cc",x"1e",x"c0"),
   238 => (x"87",x"e5",x"fd",x"49"),
   239 => (x"4b",x"70",x"86",x"c4"),
   240 => (x"c2",x"48",x"d0",x"ff"),
   241 => (x"f5",x"48",x"73",x"78"),
   242 => (x"5e",x"0e",x"87",x"c4"),
   243 => (x"0e",x"5d",x"5c",x"5b"),
   244 => (x"ff",x"c0",x"1e",x"c0"),
   245 => (x"49",x"c9",x"c1",x"f0"),
   246 => (x"d2",x"87",x"f7",x"f4"),
   247 => (x"f8",x"cc",x"c2",x"1e"),
   248 => (x"87",x"fd",x"fc",x"49"),
   249 => (x"4c",x"c0",x"86",x"c8"),
   250 => (x"b7",x"d2",x"84",x"c1"),
   251 => (x"87",x"f8",x"04",x"ac"),
   252 => (x"97",x"f8",x"cc",x"c2"),
   253 => (x"c0",x"c3",x"49",x"bf"),
   254 => (x"a9",x"c0",x"c1",x"99"),
   255 => (x"87",x"e7",x"c0",x"05"),
   256 => (x"97",x"ff",x"cc",x"c2"),
   257 => (x"31",x"d0",x"49",x"bf"),
   258 => (x"97",x"c0",x"cd",x"c2"),
   259 => (x"32",x"c8",x"4a",x"bf"),
   260 => (x"cd",x"c2",x"b1",x"72"),
   261 => (x"4a",x"bf",x"97",x"c1"),
   262 => (x"cf",x"4c",x"71",x"b1"),
   263 => (x"9c",x"ff",x"ff",x"ff"),
   264 => (x"34",x"ca",x"84",x"c1"),
   265 => (x"c2",x"87",x"e7",x"c1"),
   266 => (x"bf",x"97",x"c1",x"cd"),
   267 => (x"c6",x"31",x"c1",x"49"),
   268 => (x"c2",x"cd",x"c2",x"99"),
   269 => (x"c7",x"4a",x"bf",x"97"),
   270 => (x"b1",x"72",x"2a",x"b7"),
   271 => (x"97",x"fd",x"cc",x"c2"),
   272 => (x"cf",x"4d",x"4a",x"bf"),
   273 => (x"fe",x"cc",x"c2",x"9d"),
   274 => (x"c3",x"4a",x"bf",x"97"),
   275 => (x"c2",x"32",x"ca",x"9a"),
   276 => (x"bf",x"97",x"ff",x"cc"),
   277 => (x"73",x"33",x"c2",x"4b"),
   278 => (x"c0",x"cd",x"c2",x"b2"),
   279 => (x"c3",x"4b",x"bf",x"97"),
   280 => (x"b7",x"c6",x"9b",x"c0"),
   281 => (x"c2",x"b2",x"73",x"2b"),
   282 => (x"71",x"48",x"c1",x"81"),
   283 => (x"c1",x"49",x"70",x"30"),
   284 => (x"70",x"30",x"75",x"48"),
   285 => (x"c1",x"4c",x"72",x"4d"),
   286 => (x"c8",x"94",x"71",x"84"),
   287 => (x"06",x"ad",x"b7",x"c0"),
   288 => (x"34",x"c1",x"87",x"cc"),
   289 => (x"c0",x"c8",x"2d",x"b7"),
   290 => (x"ff",x"01",x"ad",x"b7"),
   291 => (x"48",x"74",x"87",x"f4"),
   292 => (x"0e",x"87",x"f7",x"f1"),
   293 => (x"5d",x"5c",x"5b",x"5e"),
   294 => (x"c2",x"86",x"f8",x"0e"),
   295 => (x"c0",x"48",x"de",x"d5"),
   296 => (x"d6",x"cd",x"c2",x"78"),
   297 => (x"fb",x"49",x"c0",x"1e"),
   298 => (x"86",x"c4",x"87",x"de"),
   299 => (x"c5",x"05",x"98",x"70"),
   300 => (x"c9",x"48",x"c0",x"87"),
   301 => (x"4d",x"c0",x"87",x"c0"),
   302 => (x"ed",x"c0",x"7e",x"c1"),
   303 => (x"c2",x"49",x"bf",x"eb"),
   304 => (x"71",x"4a",x"cc",x"ce"),
   305 => (x"e0",x"ee",x"4b",x"c8"),
   306 => (x"05",x"98",x"70",x"87"),
   307 => (x"7e",x"c0",x"87",x"c2"),
   308 => (x"bf",x"e7",x"ed",x"c0"),
   309 => (x"e8",x"ce",x"c2",x"49"),
   310 => (x"4b",x"c8",x"71",x"4a"),
   311 => (x"70",x"87",x"ca",x"ee"),
   312 => (x"87",x"c2",x"05",x"98"),
   313 => (x"02",x"6e",x"7e",x"c0"),
   314 => (x"c2",x"87",x"fd",x"c0"),
   315 => (x"4d",x"bf",x"dc",x"d4"),
   316 => (x"9f",x"d4",x"d5",x"c2"),
   317 => (x"c5",x"48",x"7e",x"bf"),
   318 => (x"05",x"a8",x"ea",x"d6"),
   319 => (x"d4",x"c2",x"87",x"c7"),
   320 => (x"ce",x"4d",x"bf",x"dc"),
   321 => (x"ca",x"48",x"6e",x"87"),
   322 => (x"02",x"a8",x"d5",x"e9"),
   323 => (x"48",x"c0",x"87",x"c5"),
   324 => (x"c2",x"87",x"e3",x"c7"),
   325 => (x"75",x"1e",x"d6",x"cd"),
   326 => (x"87",x"ec",x"f9",x"49"),
   327 => (x"98",x"70",x"86",x"c4"),
   328 => (x"c0",x"87",x"c5",x"05"),
   329 => (x"87",x"ce",x"c7",x"48"),
   330 => (x"bf",x"e7",x"ed",x"c0"),
   331 => (x"e8",x"ce",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f2",x"ec"),
   334 => (x"87",x"c8",x"05",x"98"),
   335 => (x"48",x"de",x"d5",x"c2"),
   336 => (x"87",x"da",x"78",x"c1"),
   337 => (x"bf",x"eb",x"ed",x"c0"),
   338 => (x"cc",x"ce",x"c2",x"49"),
   339 => (x"4b",x"c8",x"71",x"4a"),
   340 => (x"70",x"87",x"d6",x"ec"),
   341 => (x"c5",x"c0",x"02",x"98"),
   342 => (x"c6",x"48",x"c0",x"87"),
   343 => (x"d5",x"c2",x"87",x"d8"),
   344 => (x"49",x"bf",x"97",x"d4"),
   345 => (x"05",x"a9",x"d5",x"c1"),
   346 => (x"c2",x"87",x"cd",x"c0"),
   347 => (x"bf",x"97",x"d5",x"d5"),
   348 => (x"a9",x"ea",x"c2",x"49"),
   349 => (x"87",x"c5",x"c0",x"02"),
   350 => (x"f9",x"c5",x"48",x"c0"),
   351 => (x"d6",x"cd",x"c2",x"87"),
   352 => (x"48",x"7e",x"bf",x"97"),
   353 => (x"02",x"a8",x"e9",x"c3"),
   354 => (x"6e",x"87",x"ce",x"c0"),
   355 => (x"a8",x"eb",x"c3",x"48"),
   356 => (x"87",x"c5",x"c0",x"02"),
   357 => (x"dd",x"c5",x"48",x"c0"),
   358 => (x"e1",x"cd",x"c2",x"87"),
   359 => (x"99",x"49",x"bf",x"97"),
   360 => (x"87",x"cc",x"c0",x"05"),
   361 => (x"97",x"e2",x"cd",x"c2"),
   362 => (x"a9",x"c2",x"49",x"bf"),
   363 => (x"87",x"c5",x"c0",x"02"),
   364 => (x"c1",x"c5",x"48",x"c0"),
   365 => (x"e3",x"cd",x"c2",x"87"),
   366 => (x"c2",x"48",x"bf",x"97"),
   367 => (x"70",x"58",x"da",x"d5"),
   368 => (x"88",x"c1",x"48",x"4c"),
   369 => (x"58",x"de",x"d5",x"c2"),
   370 => (x"97",x"e4",x"cd",x"c2"),
   371 => (x"81",x"75",x"49",x"bf"),
   372 => (x"97",x"e5",x"cd",x"c2"),
   373 => (x"32",x"c8",x"4a",x"bf"),
   374 => (x"c2",x"7e",x"a1",x"72"),
   375 => (x"6e",x"48",x"eb",x"d9"),
   376 => (x"e6",x"cd",x"c2",x"78"),
   377 => (x"c8",x"48",x"bf",x"97"),
   378 => (x"d5",x"c2",x"58",x"a6"),
   379 => (x"c2",x"02",x"bf",x"de"),
   380 => (x"ed",x"c0",x"87",x"cf"),
   381 => (x"c2",x"49",x"bf",x"e7"),
   382 => (x"71",x"4a",x"e8",x"ce"),
   383 => (x"e8",x"e9",x"4b",x"c8"),
   384 => (x"02",x"98",x"70",x"87"),
   385 => (x"c0",x"87",x"c5",x"c0"),
   386 => (x"87",x"ea",x"c3",x"48"),
   387 => (x"bf",x"d6",x"d5",x"c2"),
   388 => (x"ff",x"d9",x"c2",x"4c"),
   389 => (x"fb",x"cd",x"c2",x"5c"),
   390 => (x"c8",x"49",x"bf",x"97"),
   391 => (x"fa",x"cd",x"c2",x"31"),
   392 => (x"a1",x"4a",x"bf",x"97"),
   393 => (x"fc",x"cd",x"c2",x"49"),
   394 => (x"d0",x"4a",x"bf",x"97"),
   395 => (x"49",x"a1",x"72",x"32"),
   396 => (x"97",x"fd",x"cd",x"c2"),
   397 => (x"32",x"d8",x"4a",x"bf"),
   398 => (x"c4",x"49",x"a1",x"72"),
   399 => (x"d9",x"c2",x"91",x"66"),
   400 => (x"c2",x"81",x"bf",x"eb"),
   401 => (x"c2",x"59",x"f3",x"d9"),
   402 => (x"bf",x"97",x"c3",x"ce"),
   403 => (x"c2",x"32",x"c8",x"4a"),
   404 => (x"bf",x"97",x"c2",x"ce"),
   405 => (x"c2",x"4a",x"a2",x"4b"),
   406 => (x"bf",x"97",x"c4",x"ce"),
   407 => (x"73",x"33",x"d0",x"4b"),
   408 => (x"ce",x"c2",x"4a",x"a2"),
   409 => (x"4b",x"bf",x"97",x"c5"),
   410 => (x"33",x"d8",x"9b",x"cf"),
   411 => (x"c2",x"4a",x"a2",x"73"),
   412 => (x"c2",x"5a",x"f7",x"d9"),
   413 => (x"c2",x"92",x"74",x"8a"),
   414 => (x"72",x"48",x"f7",x"d9"),
   415 => (x"c1",x"c1",x"78",x"a1"),
   416 => (x"e8",x"cd",x"c2",x"87"),
   417 => (x"c8",x"49",x"bf",x"97"),
   418 => (x"e7",x"cd",x"c2",x"31"),
   419 => (x"a1",x"4a",x"bf",x"97"),
   420 => (x"c7",x"31",x"c5",x"49"),
   421 => (x"29",x"c9",x"81",x"ff"),
   422 => (x"59",x"ff",x"d9",x"c2"),
   423 => (x"97",x"ed",x"cd",x"c2"),
   424 => (x"32",x"c8",x"4a",x"bf"),
   425 => (x"97",x"ec",x"cd",x"c2"),
   426 => (x"4a",x"a2",x"4b",x"bf"),
   427 => (x"6e",x"92",x"66",x"c4"),
   428 => (x"fb",x"d9",x"c2",x"82"),
   429 => (x"f3",x"d9",x"c2",x"5a"),
   430 => (x"c2",x"78",x"c0",x"48"),
   431 => (x"72",x"48",x"ef",x"d9"),
   432 => (x"d9",x"c2",x"78",x"a1"),
   433 => (x"d9",x"c2",x"48",x"ff"),
   434 => (x"c2",x"78",x"bf",x"f3"),
   435 => (x"c2",x"48",x"c3",x"da"),
   436 => (x"78",x"bf",x"f7",x"d9"),
   437 => (x"bf",x"de",x"d5",x"c2"),
   438 => (x"87",x"c9",x"c0",x"02"),
   439 => (x"30",x"c4",x"48",x"74"),
   440 => (x"c9",x"c0",x"7e",x"70"),
   441 => (x"fb",x"d9",x"c2",x"87"),
   442 => (x"30",x"c4",x"48",x"bf"),
   443 => (x"d5",x"c2",x"7e",x"70"),
   444 => (x"78",x"6e",x"48",x"e2"),
   445 => (x"8e",x"f8",x"48",x"c1"),
   446 => (x"4c",x"26",x"4d",x"26"),
   447 => (x"4f",x"26",x"4b",x"26"),
   448 => (x"5c",x"5b",x"5e",x"0e"),
   449 => (x"4a",x"71",x"0e",x"5d"),
   450 => (x"bf",x"de",x"d5",x"c2"),
   451 => (x"72",x"87",x"cb",x"02"),
   452 => (x"72",x"2b",x"c7",x"4b"),
   453 => (x"9d",x"ff",x"c1",x"4d"),
   454 => (x"4b",x"72",x"87",x"c9"),
   455 => (x"4d",x"72",x"2b",x"c8"),
   456 => (x"c2",x"9d",x"ff",x"c3"),
   457 => (x"83",x"bf",x"eb",x"d9"),
   458 => (x"bf",x"e3",x"ed",x"c0"),
   459 => (x"87",x"d9",x"02",x"ab"),
   460 => (x"5b",x"e7",x"ed",x"c0"),
   461 => (x"1e",x"d6",x"cd",x"c2"),
   462 => (x"cb",x"f1",x"49",x"73"),
   463 => (x"70",x"86",x"c4",x"87"),
   464 => (x"87",x"c5",x"05",x"98"),
   465 => (x"e6",x"c0",x"48",x"c0"),
   466 => (x"de",x"d5",x"c2",x"87"),
   467 => (x"87",x"d2",x"02",x"bf"),
   468 => (x"91",x"c4",x"49",x"75"),
   469 => (x"81",x"d6",x"cd",x"c2"),
   470 => (x"ff",x"cf",x"4c",x"69"),
   471 => (x"9c",x"ff",x"ff",x"ff"),
   472 => (x"49",x"75",x"87",x"cb"),
   473 => (x"cd",x"c2",x"91",x"c2"),
   474 => (x"69",x"9f",x"81",x"d6"),
   475 => (x"fe",x"48",x"74",x"4c"),
   476 => (x"5e",x"0e",x"87",x"c6"),
   477 => (x"0e",x"5d",x"5c",x"5b"),
   478 => (x"4c",x"71",x"86",x"f8"),
   479 => (x"87",x"c5",x"05",x"9c"),
   480 => (x"c1",x"c3",x"48",x"c0"),
   481 => (x"7e",x"a4",x"c8",x"87"),
   482 => (x"d8",x"78",x"c0",x"48"),
   483 => (x"87",x"c7",x"02",x"66"),
   484 => (x"bf",x"97",x"66",x"d8"),
   485 => (x"c0",x"87",x"c5",x"05"),
   486 => (x"87",x"ea",x"c2",x"48"),
   487 => (x"49",x"c1",x"1e",x"c0"),
   488 => (x"87",x"e6",x"c7",x"49"),
   489 => (x"4d",x"70",x"86",x"c4"),
   490 => (x"c2",x"c1",x"02",x"9d"),
   491 => (x"e6",x"d5",x"c2",x"87"),
   492 => (x"49",x"66",x"d8",x"4a"),
   493 => (x"70",x"87",x"d7",x"e2"),
   494 => (x"f2",x"c0",x"02",x"98"),
   495 => (x"d8",x"4a",x"75",x"87"),
   496 => (x"4b",x"cb",x"49",x"66"),
   497 => (x"70",x"87",x"fc",x"e2"),
   498 => (x"e2",x"c0",x"02",x"98"),
   499 => (x"75",x"1e",x"c0",x"87"),
   500 => (x"87",x"c7",x"02",x"9d"),
   501 => (x"c0",x"48",x"a6",x"c8"),
   502 => (x"c8",x"87",x"c5",x"78"),
   503 => (x"78",x"c1",x"48",x"a6"),
   504 => (x"c6",x"49",x"66",x"c8"),
   505 => (x"86",x"c4",x"87",x"e4"),
   506 => (x"05",x"9d",x"4d",x"70"),
   507 => (x"75",x"87",x"fe",x"fe"),
   508 => (x"cf",x"c1",x"02",x"9d"),
   509 => (x"49",x"a5",x"dc",x"87"),
   510 => (x"78",x"69",x"48",x"6e"),
   511 => (x"c4",x"49",x"a5",x"da"),
   512 => (x"a4",x"c4",x"48",x"a6"),
   513 => (x"48",x"69",x"9f",x"78"),
   514 => (x"78",x"08",x"66",x"c4"),
   515 => (x"bf",x"de",x"d5",x"c2"),
   516 => (x"d4",x"87",x"d2",x"02"),
   517 => (x"69",x"9f",x"49",x"a5"),
   518 => (x"ff",x"ff",x"c0",x"49"),
   519 => (x"d0",x"48",x"71",x"99"),
   520 => (x"c2",x"7e",x"70",x"30"),
   521 => (x"6e",x"7e",x"c0",x"87"),
   522 => (x"66",x"c4",x"48",x"49"),
   523 => (x"66",x"c4",x"80",x"bf"),
   524 => (x"7c",x"c0",x"78",x"08"),
   525 => (x"c4",x"49",x"a4",x"cc"),
   526 => (x"d0",x"79",x"bf",x"66"),
   527 => (x"79",x"c0",x"49",x"a4"),
   528 => (x"87",x"c2",x"48",x"c1"),
   529 => (x"8e",x"f8",x"48",x"c0"),
   530 => (x"0e",x"87",x"ed",x"fa"),
   531 => (x"5d",x"5c",x"5b",x"5e"),
   532 => (x"9c",x"4c",x"71",x"0e"),
   533 => (x"87",x"cb",x"c1",x"02"),
   534 => (x"69",x"49",x"a4",x"c8"),
   535 => (x"87",x"c3",x"c1",x"02"),
   536 => (x"6c",x"4a",x"66",x"d0"),
   537 => (x"48",x"a6",x"d0",x"49"),
   538 => (x"4d",x"78",x"a1",x"72"),
   539 => (x"da",x"d5",x"c2",x"b9"),
   540 => (x"ba",x"ff",x"4a",x"bf"),
   541 => (x"99",x"71",x"99",x"72"),
   542 => (x"87",x"e4",x"c0",x"02"),
   543 => (x"6b",x"4b",x"a4",x"c4"),
   544 => (x"87",x"fc",x"f9",x"49"),
   545 => (x"d5",x"c2",x"7b",x"70"),
   546 => (x"6c",x"49",x"bf",x"d6"),
   547 => (x"75",x"7c",x"71",x"81"),
   548 => (x"da",x"d5",x"c2",x"b9"),
   549 => (x"ba",x"ff",x"4a",x"bf"),
   550 => (x"99",x"71",x"99",x"72"),
   551 => (x"87",x"dc",x"ff",x"05"),
   552 => (x"f9",x"7c",x"66",x"d0"),
   553 => (x"73",x"1e",x"87",x"d2"),
   554 => (x"9b",x"4b",x"71",x"1e"),
   555 => (x"c8",x"87",x"c7",x"02"),
   556 => (x"05",x"69",x"49",x"a3"),
   557 => (x"48",x"c0",x"87",x"c5"),
   558 => (x"c2",x"87",x"f6",x"c0"),
   559 => (x"49",x"bf",x"ef",x"d9"),
   560 => (x"6a",x"4a",x"a3",x"c4"),
   561 => (x"c2",x"8a",x"c2",x"4a"),
   562 => (x"92",x"bf",x"d6",x"d5"),
   563 => (x"c2",x"49",x"a1",x"72"),
   564 => (x"4a",x"bf",x"da",x"d5"),
   565 => (x"a1",x"72",x"9a",x"6b"),
   566 => (x"e7",x"ed",x"c0",x"49"),
   567 => (x"1e",x"66",x"c8",x"59"),
   568 => (x"87",x"e4",x"ea",x"71"),
   569 => (x"98",x"70",x"86",x"c4"),
   570 => (x"c0",x"87",x"c4",x"05"),
   571 => (x"c1",x"87",x"c2",x"48"),
   572 => (x"87",x"c8",x"f8",x"48"),
   573 => (x"71",x"1e",x"73",x"1e"),
   574 => (x"c0",x"02",x"9b",x"4b"),
   575 => (x"da",x"c2",x"87",x"e4"),
   576 => (x"4a",x"73",x"5b",x"c3"),
   577 => (x"d5",x"c2",x"8a",x"c2"),
   578 => (x"92",x"49",x"bf",x"d6"),
   579 => (x"bf",x"ef",x"d9",x"c2"),
   580 => (x"c2",x"80",x"72",x"48"),
   581 => (x"71",x"58",x"c7",x"da"),
   582 => (x"c2",x"30",x"c4",x"48"),
   583 => (x"c0",x"58",x"e6",x"d5"),
   584 => (x"d9",x"c2",x"87",x"ed"),
   585 => (x"d9",x"c2",x"48",x"ff"),
   586 => (x"c2",x"78",x"bf",x"f3"),
   587 => (x"c2",x"48",x"c3",x"da"),
   588 => (x"78",x"bf",x"f7",x"d9"),
   589 => (x"bf",x"de",x"d5",x"c2"),
   590 => (x"c2",x"87",x"c9",x"02"),
   591 => (x"49",x"bf",x"d6",x"d5"),
   592 => (x"87",x"c7",x"31",x"c4"),
   593 => (x"bf",x"fb",x"d9",x"c2"),
   594 => (x"c2",x"31",x"c4",x"49"),
   595 => (x"f6",x"59",x"e6",x"d5"),
   596 => (x"5e",x"0e",x"87",x"ea"),
   597 => (x"71",x"0e",x"5c",x"5b"),
   598 => (x"72",x"4b",x"c0",x"4a"),
   599 => (x"e1",x"c0",x"02",x"9a"),
   600 => (x"49",x"a2",x"da",x"87"),
   601 => (x"c2",x"4b",x"69",x"9f"),
   602 => (x"02",x"bf",x"de",x"d5"),
   603 => (x"a2",x"d4",x"87",x"cf"),
   604 => (x"49",x"69",x"9f",x"49"),
   605 => (x"ff",x"ff",x"c0",x"4c"),
   606 => (x"c2",x"34",x"d0",x"9c"),
   607 => (x"74",x"4c",x"c0",x"87"),
   608 => (x"49",x"73",x"b3",x"49"),
   609 => (x"f5",x"87",x"ed",x"fd"),
   610 => (x"5e",x"0e",x"87",x"f0"),
   611 => (x"0e",x"5d",x"5c",x"5b"),
   612 => (x"4a",x"71",x"86",x"f4"),
   613 => (x"9a",x"72",x"7e",x"c0"),
   614 => (x"c2",x"87",x"d8",x"02"),
   615 => (x"c0",x"48",x"d2",x"cd"),
   616 => (x"ca",x"cd",x"c2",x"78"),
   617 => (x"c3",x"da",x"c2",x"48"),
   618 => (x"cd",x"c2",x"78",x"bf"),
   619 => (x"d9",x"c2",x"48",x"ce"),
   620 => (x"c2",x"78",x"bf",x"ff"),
   621 => (x"c0",x"48",x"f3",x"d5"),
   622 => (x"e2",x"d5",x"c2",x"50"),
   623 => (x"cd",x"c2",x"49",x"bf"),
   624 => (x"71",x"4a",x"bf",x"d2"),
   625 => (x"c9",x"c4",x"03",x"aa"),
   626 => (x"cf",x"49",x"72",x"87"),
   627 => (x"e9",x"c0",x"05",x"99"),
   628 => (x"e3",x"ed",x"c0",x"87"),
   629 => (x"ca",x"cd",x"c2",x"48"),
   630 => (x"cd",x"c2",x"78",x"bf"),
   631 => (x"cd",x"c2",x"1e",x"d6"),
   632 => (x"c2",x"49",x"bf",x"ca"),
   633 => (x"c1",x"48",x"ca",x"cd"),
   634 => (x"e6",x"71",x"78",x"a1"),
   635 => (x"86",x"c4",x"87",x"da"),
   636 => (x"48",x"df",x"ed",x"c0"),
   637 => (x"78",x"d6",x"cd",x"c2"),
   638 => (x"ed",x"c0",x"87",x"cc"),
   639 => (x"c0",x"48",x"bf",x"df"),
   640 => (x"ed",x"c0",x"80",x"e0"),
   641 => (x"cd",x"c2",x"58",x"e3"),
   642 => (x"c1",x"48",x"bf",x"d2"),
   643 => (x"d6",x"cd",x"c2",x"80"),
   644 => (x"0b",x"5f",x"27",x"58"),
   645 => (x"97",x"bf",x"00",x"00"),
   646 => (x"02",x"9d",x"4d",x"bf"),
   647 => (x"c3",x"87",x"e3",x"c2"),
   648 => (x"c2",x"02",x"ad",x"e5"),
   649 => (x"ed",x"c0",x"87",x"dc"),
   650 => (x"cb",x"4b",x"bf",x"df"),
   651 => (x"4c",x"11",x"49",x"a3"),
   652 => (x"c1",x"05",x"ac",x"cf"),
   653 => (x"49",x"75",x"87",x"d2"),
   654 => (x"89",x"c1",x"99",x"df"),
   655 => (x"d5",x"c2",x"91",x"cd"),
   656 => (x"a3",x"c1",x"81",x"e6"),
   657 => (x"c3",x"51",x"12",x"4a"),
   658 => (x"51",x"12",x"4a",x"a3"),
   659 => (x"12",x"4a",x"a3",x"c5"),
   660 => (x"4a",x"a3",x"c7",x"51"),
   661 => (x"a3",x"c9",x"51",x"12"),
   662 => (x"ce",x"51",x"12",x"4a"),
   663 => (x"51",x"12",x"4a",x"a3"),
   664 => (x"12",x"4a",x"a3",x"d0"),
   665 => (x"4a",x"a3",x"d2",x"51"),
   666 => (x"a3",x"d4",x"51",x"12"),
   667 => (x"d6",x"51",x"12",x"4a"),
   668 => (x"51",x"12",x"4a",x"a3"),
   669 => (x"12",x"4a",x"a3",x"d8"),
   670 => (x"4a",x"a3",x"dc",x"51"),
   671 => (x"a3",x"de",x"51",x"12"),
   672 => (x"c1",x"51",x"12",x"4a"),
   673 => (x"87",x"fa",x"c0",x"7e"),
   674 => (x"99",x"c8",x"49",x"74"),
   675 => (x"87",x"eb",x"c0",x"05"),
   676 => (x"99",x"d0",x"49",x"74"),
   677 => (x"dc",x"87",x"d1",x"05"),
   678 => (x"cb",x"c0",x"02",x"66"),
   679 => (x"dc",x"49",x"73",x"87"),
   680 => (x"98",x"70",x"0f",x"66"),
   681 => (x"87",x"d3",x"c0",x"02"),
   682 => (x"c6",x"c0",x"05",x"6e"),
   683 => (x"e6",x"d5",x"c2",x"87"),
   684 => (x"c0",x"50",x"c0",x"48"),
   685 => (x"48",x"bf",x"df",x"ed"),
   686 => (x"c2",x"87",x"df",x"c2"),
   687 => (x"c0",x"48",x"f3",x"d5"),
   688 => (x"d5",x"c2",x"7e",x"50"),
   689 => (x"c2",x"49",x"bf",x"e2"),
   690 => (x"4a",x"bf",x"d2",x"cd"),
   691 => (x"fb",x"04",x"aa",x"71"),
   692 => (x"da",x"c2",x"87",x"f7"),
   693 => (x"c0",x"05",x"bf",x"c3"),
   694 => (x"d5",x"c2",x"87",x"c8"),
   695 => (x"c1",x"02",x"bf",x"de"),
   696 => (x"cd",x"c2",x"87",x"f6"),
   697 => (x"f0",x"49",x"bf",x"ce"),
   698 => (x"cd",x"c2",x"87",x"d6"),
   699 => (x"a6",x"c4",x"58",x"d2"),
   700 => (x"ce",x"cd",x"c2",x"48"),
   701 => (x"d5",x"c2",x"78",x"bf"),
   702 => (x"c0",x"02",x"bf",x"de"),
   703 => (x"66",x"c4",x"87",x"d8"),
   704 => (x"ff",x"ff",x"cf",x"49"),
   705 => (x"a9",x"99",x"f8",x"ff"),
   706 => (x"87",x"c5",x"c0",x"02"),
   707 => (x"e1",x"c0",x"4c",x"c0"),
   708 => (x"c0",x"4c",x"c1",x"87"),
   709 => (x"66",x"c4",x"87",x"dc"),
   710 => (x"f8",x"ff",x"cf",x"49"),
   711 => (x"c0",x"02",x"a9",x"99"),
   712 => (x"a6",x"c8",x"87",x"c8"),
   713 => (x"c0",x"78",x"c0",x"48"),
   714 => (x"a6",x"c8",x"87",x"c5"),
   715 => (x"c8",x"78",x"c1",x"48"),
   716 => (x"9c",x"74",x"4c",x"66"),
   717 => (x"87",x"e0",x"c0",x"05"),
   718 => (x"c2",x"49",x"66",x"c4"),
   719 => (x"d6",x"d5",x"c2",x"89"),
   720 => (x"c2",x"91",x"4a",x"bf"),
   721 => (x"4a",x"bf",x"ef",x"d9"),
   722 => (x"48",x"ca",x"cd",x"c2"),
   723 => (x"c2",x"78",x"a1",x"72"),
   724 => (x"c0",x"48",x"d2",x"cd"),
   725 => (x"87",x"e1",x"f9",x"78"),
   726 => (x"8e",x"f4",x"48",x"c0"),
   727 => (x"00",x"87",x"d9",x"ee"),
   728 => (x"ff",x"00",x"00",x"00"),
   729 => (x"6f",x"ff",x"ff",x"ff"),
   730 => (x"78",x"00",x"00",x"0b"),
   731 => (x"46",x"00",x"00",x"0b"),
   732 => (x"32",x"33",x"54",x"41"),
   733 => (x"00",x"20",x"20",x"20"),
   734 => (x"31",x"54",x"41",x"46"),
   735 => (x"20",x"20",x"20",x"36"),
   736 => (x"d4",x"ff",x"1e",x"00"),
   737 => (x"78",x"ff",x"c3",x"48"),
   738 => (x"4f",x"26",x"48",x"68"),
   739 => (x"48",x"d4",x"ff",x"1e"),
   740 => (x"ff",x"78",x"ff",x"c3"),
   741 => (x"e1",x"c0",x"48",x"d0"),
   742 => (x"48",x"d4",x"ff",x"78"),
   743 => (x"da",x"c2",x"78",x"d4"),
   744 => (x"d4",x"ff",x"48",x"c7"),
   745 => (x"4f",x"26",x"50",x"bf"),
   746 => (x"48",x"d0",x"ff",x"1e"),
   747 => (x"26",x"78",x"e0",x"c0"),
   748 => (x"cc",x"ff",x"1e",x"4f"),
   749 => (x"99",x"49",x"70",x"87"),
   750 => (x"c0",x"87",x"c6",x"02"),
   751 => (x"f1",x"05",x"a9",x"fb"),
   752 => (x"26",x"48",x"71",x"87"),
   753 => (x"5b",x"5e",x"0e",x"4f"),
   754 => (x"4b",x"71",x"0e",x"5c"),
   755 => (x"f0",x"fe",x"4c",x"c0"),
   756 => (x"99",x"49",x"70",x"87"),
   757 => (x"87",x"f9",x"c0",x"02"),
   758 => (x"02",x"a9",x"ec",x"c0"),
   759 => (x"c0",x"87",x"f2",x"c0"),
   760 => (x"c0",x"02",x"a9",x"fb"),
   761 => (x"66",x"cc",x"87",x"eb"),
   762 => (x"c7",x"03",x"ac",x"b7"),
   763 => (x"02",x"66",x"d0",x"87"),
   764 => (x"53",x"71",x"87",x"c2"),
   765 => (x"c2",x"02",x"99",x"71"),
   766 => (x"fe",x"84",x"c1",x"87"),
   767 => (x"49",x"70",x"87",x"c3"),
   768 => (x"87",x"cd",x"02",x"99"),
   769 => (x"02",x"a9",x"ec",x"c0"),
   770 => (x"fb",x"c0",x"87",x"c7"),
   771 => (x"d5",x"ff",x"05",x"a9"),
   772 => (x"02",x"66",x"d0",x"87"),
   773 => (x"97",x"c0",x"87",x"c3"),
   774 => (x"a9",x"ec",x"c0",x"7b"),
   775 => (x"74",x"87",x"c4",x"05"),
   776 => (x"74",x"87",x"c5",x"4a"),
   777 => (x"8a",x"0a",x"c0",x"4a"),
   778 => (x"87",x"c2",x"48",x"72"),
   779 => (x"4c",x"26",x"4d",x"26"),
   780 => (x"4f",x"26",x"4b",x"26"),
   781 => (x"87",x"c9",x"fd",x"1e"),
   782 => (x"f0",x"c0",x"4a",x"70"),
   783 => (x"87",x"c9",x"04",x"aa"),
   784 => (x"01",x"aa",x"f9",x"c0"),
   785 => (x"f0",x"c0",x"87",x"c3"),
   786 => (x"aa",x"c1",x"c1",x"8a"),
   787 => (x"c1",x"87",x"c9",x"04"),
   788 => (x"c3",x"01",x"aa",x"da"),
   789 => (x"8a",x"f7",x"c0",x"87"),
   790 => (x"4f",x"26",x"48",x"72"),
   791 => (x"5c",x"5b",x"5e",x"0e"),
   792 => (x"86",x"f8",x"0e",x"5d"),
   793 => (x"4d",x"c0",x"4c",x"71"),
   794 => (x"c0",x"87",x"e1",x"fc"),
   795 => (x"fb",x"f3",x"c0",x"4b"),
   796 => (x"c0",x"49",x"bf",x"97"),
   797 => (x"87",x"cf",x"04",x"a9"),
   798 => (x"c1",x"87",x"f6",x"fc"),
   799 => (x"fb",x"f3",x"c0",x"83"),
   800 => (x"ab",x"49",x"bf",x"97"),
   801 => (x"c0",x"87",x"f1",x"06"),
   802 => (x"bf",x"97",x"fb",x"f3"),
   803 => (x"fb",x"87",x"cf",x"02"),
   804 => (x"49",x"70",x"87",x"ef"),
   805 => (x"87",x"c6",x"02",x"99"),
   806 => (x"05",x"a9",x"ec",x"c0"),
   807 => (x"4b",x"c0",x"87",x"f1"),
   808 => (x"70",x"87",x"de",x"fb"),
   809 => (x"87",x"d9",x"fb",x"7e"),
   810 => (x"fb",x"58",x"a6",x"c8"),
   811 => (x"4a",x"70",x"87",x"d3"),
   812 => (x"a4",x"c8",x"83",x"c1"),
   813 => (x"49",x"69",x"97",x"49"),
   814 => (x"da",x"05",x"a9",x"6e"),
   815 => (x"49",x"a4",x"c9",x"87"),
   816 => (x"c4",x"49",x"69",x"97"),
   817 => (x"ce",x"05",x"a9",x"66"),
   818 => (x"49",x"a4",x"ca",x"87"),
   819 => (x"aa",x"49",x"69",x"97"),
   820 => (x"c1",x"87",x"c4",x"05"),
   821 => (x"6e",x"87",x"d4",x"4d"),
   822 => (x"a8",x"ec",x"c0",x"48"),
   823 => (x"6e",x"87",x"c8",x"02"),
   824 => (x"a8",x"fb",x"c0",x"48"),
   825 => (x"c0",x"87",x"c4",x"05"),
   826 => (x"75",x"4d",x"c1",x"4b"),
   827 => (x"ef",x"fe",x"02",x"9d"),
   828 => (x"87",x"f4",x"fa",x"87"),
   829 => (x"8e",x"f8",x"48",x"73"),
   830 => (x"00",x"87",x"f1",x"fc"),
   831 => (x"5c",x"5b",x"5e",x"0e"),
   832 => (x"86",x"f8",x"0e",x"5d"),
   833 => (x"d4",x"ff",x"7e",x"71"),
   834 => (x"c2",x"1e",x"6e",x"4b"),
   835 => (x"e9",x"49",x"cc",x"da"),
   836 => (x"86",x"c4",x"87",x"e0"),
   837 => (x"c4",x"02",x"98",x"70"),
   838 => (x"dd",x"c1",x"87",x"ea"),
   839 => (x"6e",x"4d",x"bf",x"e2"),
   840 => (x"87",x"f8",x"fc",x"49"),
   841 => (x"70",x"58",x"a6",x"c8"),
   842 => (x"87",x"c5",x"05",x"98"),
   843 => (x"c1",x"48",x"a6",x"c4"),
   844 => (x"48",x"d0",x"ff",x"78"),
   845 => (x"d5",x"c1",x"78",x"c5"),
   846 => (x"49",x"66",x"c4",x"7b"),
   847 => (x"31",x"c6",x"89",x"c1"),
   848 => (x"97",x"e0",x"dd",x"c1"),
   849 => (x"71",x"48",x"4a",x"bf"),
   850 => (x"ff",x"7b",x"70",x"b0"),
   851 => (x"78",x"c4",x"48",x"d0"),
   852 => (x"97",x"c7",x"da",x"c2"),
   853 => (x"99",x"d0",x"49",x"bf"),
   854 => (x"c5",x"87",x"d7",x"02"),
   855 => (x"7b",x"d6",x"c1",x"78"),
   856 => (x"ff",x"c3",x"4a",x"c0"),
   857 => (x"c0",x"82",x"c1",x"7b"),
   858 => (x"f5",x"04",x"aa",x"e0"),
   859 => (x"48",x"d0",x"ff",x"87"),
   860 => (x"ff",x"c3",x"78",x"c4"),
   861 => (x"48",x"d0",x"ff",x"7b"),
   862 => (x"d3",x"c1",x"78",x"c5"),
   863 => (x"c4",x"7b",x"c1",x"7b"),
   864 => (x"ad",x"b7",x"c0",x"78"),
   865 => (x"87",x"eb",x"c2",x"06"),
   866 => (x"bf",x"d4",x"da",x"c2"),
   867 => (x"02",x"9c",x"8d",x"4c"),
   868 => (x"c2",x"87",x"c2",x"c2"),
   869 => (x"c4",x"7e",x"d6",x"cd"),
   870 => (x"c0",x"c8",x"48",x"a6"),
   871 => (x"b7",x"c0",x"8c",x"78"),
   872 => (x"87",x"c6",x"03",x"ac"),
   873 => (x"78",x"a4",x"c0",x"c8"),
   874 => (x"da",x"c2",x"4c",x"c0"),
   875 => (x"49",x"bf",x"97",x"c7"),
   876 => (x"d0",x"02",x"99",x"d0"),
   877 => (x"c2",x"1e",x"c0",x"87"),
   878 => (x"eb",x"49",x"cc",x"da"),
   879 => (x"86",x"c4",x"87",x"e8"),
   880 => (x"f5",x"c0",x"4a",x"70"),
   881 => (x"d6",x"cd",x"c2",x"87"),
   882 => (x"cc",x"da",x"c2",x"1e"),
   883 => (x"87",x"d6",x"eb",x"49"),
   884 => (x"4a",x"70",x"86",x"c4"),
   885 => (x"c8",x"48",x"d0",x"ff"),
   886 => (x"d4",x"c1",x"78",x"c5"),
   887 => (x"bf",x"97",x"6e",x"7b"),
   888 => (x"c1",x"48",x"6e",x"7b"),
   889 => (x"c4",x"7e",x"70",x"80"),
   890 => (x"88",x"c1",x"48",x"66"),
   891 => (x"70",x"58",x"a6",x"c8"),
   892 => (x"e8",x"ff",x"05",x"98"),
   893 => (x"48",x"d0",x"ff",x"87"),
   894 => (x"9a",x"72",x"78",x"c4"),
   895 => (x"c0",x"87",x"c5",x"05"),
   896 => (x"87",x"c2",x"c1",x"48"),
   897 => (x"da",x"c2",x"1e",x"c1"),
   898 => (x"fe",x"e8",x"49",x"cc"),
   899 => (x"74",x"86",x"c4",x"87"),
   900 => (x"fe",x"fd",x"05",x"9c"),
   901 => (x"ad",x"b7",x"c0",x"87"),
   902 => (x"c2",x"87",x"d1",x"06"),
   903 => (x"c0",x"48",x"cc",x"da"),
   904 => (x"c0",x"80",x"d0",x"78"),
   905 => (x"c2",x"80",x"f4",x"78"),
   906 => (x"78",x"bf",x"d8",x"da"),
   907 => (x"01",x"ad",x"b7",x"c0"),
   908 => (x"ff",x"87",x"d5",x"fd"),
   909 => (x"78",x"c5",x"48",x"d0"),
   910 => (x"c0",x"7b",x"d3",x"c1"),
   911 => (x"c1",x"78",x"c4",x"7b"),
   912 => (x"87",x"c2",x"c0",x"48"),
   913 => (x"8e",x"f8",x"48",x"c0"),
   914 => (x"4c",x"26",x"4d",x"26"),
   915 => (x"4f",x"26",x"4b",x"26"),
   916 => (x"5c",x"5b",x"5e",x"0e"),
   917 => (x"71",x"1e",x"0e",x"5d"),
   918 => (x"4d",x"4c",x"c0",x"4b"),
   919 => (x"e8",x"c0",x"04",x"ab"),
   920 => (x"dc",x"f1",x"c0",x"87"),
   921 => (x"02",x"9d",x"75",x"1e"),
   922 => (x"4a",x"c0",x"87",x"c4"),
   923 => (x"4a",x"c1",x"87",x"c2"),
   924 => (x"d5",x"ec",x"49",x"72"),
   925 => (x"70",x"86",x"c4",x"87"),
   926 => (x"6e",x"84",x"c1",x"7e"),
   927 => (x"73",x"87",x"c2",x"05"),
   928 => (x"73",x"85",x"c1",x"4c"),
   929 => (x"d8",x"ff",x"06",x"ac"),
   930 => (x"26",x"48",x"6e",x"87"),
   931 => (x"1e",x"87",x"f9",x"fe"),
   932 => (x"66",x"c4",x"4a",x"71"),
   933 => (x"72",x"87",x"c5",x"05"),
   934 => (x"87",x"e0",x"f9",x"49"),
   935 => (x"5e",x"0e",x"4f",x"26"),
   936 => (x"0e",x"5d",x"5c",x"5b"),
   937 => (x"49",x"4c",x"71",x"1e"),
   938 => (x"da",x"c2",x"91",x"de"),
   939 => (x"85",x"71",x"4d",x"f4"),
   940 => (x"c1",x"02",x"6d",x"97"),
   941 => (x"da",x"c2",x"87",x"dc"),
   942 => (x"74",x"49",x"bf",x"e0"),
   943 => (x"cf",x"fe",x"71",x"81"),
   944 => (x"48",x"7e",x"70",x"87"),
   945 => (x"f2",x"c0",x"02",x"98"),
   946 => (x"e8",x"da",x"c2",x"87"),
   947 => (x"cb",x"4a",x"70",x"4b"),
   948 => (x"d2",x"c7",x"ff",x"49"),
   949 => (x"cb",x"4b",x"74",x"87"),
   950 => (x"f4",x"dd",x"c1",x"93"),
   951 => (x"c0",x"83",x"c4",x"83"),
   952 => (x"74",x"7b",x"d6",x"fc"),
   953 => (x"ec",x"c0",x"c1",x"49"),
   954 => (x"c1",x"7b",x"75",x"87"),
   955 => (x"bf",x"97",x"e1",x"dd"),
   956 => (x"da",x"c2",x"1e",x"49"),
   957 => (x"d6",x"fe",x"49",x"e8"),
   958 => (x"74",x"86",x"c4",x"87"),
   959 => (x"d4",x"c0",x"c1",x"49"),
   960 => (x"c1",x"49",x"c0",x"87"),
   961 => (x"c2",x"87",x"f3",x"c1"),
   962 => (x"c0",x"48",x"c8",x"da"),
   963 => (x"dd",x"49",x"c1",x"78"),
   964 => (x"fc",x"26",x"87",x"f9"),
   965 => (x"6f",x"4c",x"87",x"f2"),
   966 => (x"6e",x"69",x"64",x"61"),
   967 => (x"2e",x"2e",x"2e",x"67"),
   968 => (x"1e",x"73",x"1e",x"00"),
   969 => (x"c2",x"49",x"4a",x"71"),
   970 => (x"81",x"bf",x"e0",x"da"),
   971 => (x"87",x"e0",x"fc",x"71"),
   972 => (x"02",x"9b",x"4b",x"70"),
   973 => (x"e8",x"49",x"87",x"c4"),
   974 => (x"da",x"c2",x"87",x"d8"),
   975 => (x"78",x"c0",x"48",x"e0"),
   976 => (x"c6",x"dd",x"49",x"c1"),
   977 => (x"87",x"c4",x"fc",x"87"),
   978 => (x"c1",x"49",x"c0",x"1e"),
   979 => (x"26",x"87",x"eb",x"c0"),
   980 => (x"4a",x"71",x"1e",x"4f"),
   981 => (x"c1",x"91",x"cb",x"49"),
   982 => (x"c8",x"81",x"f4",x"dd"),
   983 => (x"c2",x"48",x"11",x"81"),
   984 => (x"c2",x"58",x"cc",x"da"),
   985 => (x"c0",x"48",x"e0",x"da"),
   986 => (x"dc",x"49",x"c1",x"78"),
   987 => (x"4f",x"26",x"87",x"dd"),
   988 => (x"02",x"99",x"71",x"1e"),
   989 => (x"df",x"c1",x"87",x"d2"),
   990 => (x"50",x"c0",x"48",x"c9"),
   991 => (x"fd",x"c0",x"80",x"f7"),
   992 => (x"dd",x"c1",x"40",x"d1"),
   993 => (x"87",x"ce",x"78",x"ed"),
   994 => (x"48",x"c5",x"df",x"c1"),
   995 => (x"78",x"e6",x"dd",x"c1"),
   996 => (x"fd",x"c0",x"80",x"fc"),
   997 => (x"4f",x"26",x"78",x"c8"),
   998 => (x"5c",x"5b",x"5e",x"0e"),
   999 => (x"86",x"f4",x"0e",x"5d"),
  1000 => (x"4d",x"d6",x"cd",x"c2"),
  1001 => (x"a6",x"c4",x"4c",x"c0"),
  1002 => (x"c2",x"78",x"c0",x"48"),
  1003 => (x"48",x"bf",x"e0",x"da"),
  1004 => (x"c1",x"06",x"a8",x"c0"),
  1005 => (x"cd",x"c2",x"87",x"c0"),
  1006 => (x"02",x"98",x"48",x"d6"),
  1007 => (x"c0",x"87",x"f7",x"c0"),
  1008 => (x"c8",x"1e",x"dc",x"f1"),
  1009 => (x"87",x"c7",x"02",x"66"),
  1010 => (x"c0",x"48",x"a6",x"c4"),
  1011 => (x"c4",x"87",x"c5",x"78"),
  1012 => (x"78",x"c1",x"48",x"a6"),
  1013 => (x"e6",x"49",x"66",x"c4"),
  1014 => (x"86",x"c4",x"87",x"f0"),
  1015 => (x"84",x"c1",x"4d",x"70"),
  1016 => (x"c1",x"48",x"66",x"c4"),
  1017 => (x"58",x"a6",x"c8",x"80"),
  1018 => (x"bf",x"e0",x"da",x"c2"),
  1019 => (x"87",x"c6",x"03",x"ac"),
  1020 => (x"ff",x"05",x"9d",x"75"),
  1021 => (x"4c",x"c0",x"87",x"c9"),
  1022 => (x"c3",x"02",x"9d",x"75"),
  1023 => (x"f1",x"c0",x"87",x"dc"),
  1024 => (x"66",x"c8",x"1e",x"dc"),
  1025 => (x"cc",x"87",x"c7",x"02"),
  1026 => (x"78",x"c0",x"48",x"a6"),
  1027 => (x"a6",x"cc",x"87",x"c5"),
  1028 => (x"cc",x"78",x"c1",x"48"),
  1029 => (x"f1",x"e5",x"49",x"66"),
  1030 => (x"70",x"86",x"c4",x"87"),
  1031 => (x"02",x"98",x"48",x"7e"),
  1032 => (x"49",x"87",x"e4",x"c2"),
  1033 => (x"69",x"97",x"81",x"cb"),
  1034 => (x"02",x"99",x"d0",x"49"),
  1035 => (x"74",x"87",x"d4",x"c1"),
  1036 => (x"c1",x"91",x"cb",x"49"),
  1037 => (x"c0",x"81",x"f4",x"dd"),
  1038 => (x"c8",x"79",x"e1",x"fc"),
  1039 => (x"51",x"ff",x"c3",x"81"),
  1040 => (x"91",x"de",x"49",x"74"),
  1041 => (x"4d",x"f4",x"da",x"c2"),
  1042 => (x"c1",x"c2",x"85",x"71"),
  1043 => (x"a5",x"c1",x"7d",x"97"),
  1044 => (x"51",x"e0",x"c0",x"49"),
  1045 => (x"97",x"e6",x"d5",x"c2"),
  1046 => (x"87",x"d2",x"02",x"bf"),
  1047 => (x"a5",x"c2",x"84",x"c1"),
  1048 => (x"e6",x"d5",x"c2",x"4b"),
  1049 => (x"ff",x"49",x"db",x"4a"),
  1050 => (x"c1",x"87",x"fc",x"c0"),
  1051 => (x"a5",x"cd",x"87",x"d9"),
  1052 => (x"c1",x"51",x"c0",x"49"),
  1053 => (x"4b",x"a5",x"c2",x"84"),
  1054 => (x"49",x"cb",x"4a",x"6e"),
  1055 => (x"87",x"e7",x"c0",x"ff"),
  1056 => (x"74",x"87",x"c4",x"c1"),
  1057 => (x"c1",x"91",x"cb",x"49"),
  1058 => (x"c0",x"81",x"f4",x"dd"),
  1059 => (x"c2",x"79",x"de",x"fa"),
  1060 => (x"bf",x"97",x"e6",x"d5"),
  1061 => (x"74",x"87",x"d8",x"02"),
  1062 => (x"c1",x"91",x"de",x"49"),
  1063 => (x"f4",x"da",x"c2",x"84"),
  1064 => (x"c2",x"83",x"71",x"4b"),
  1065 => (x"dd",x"4a",x"e6",x"d5"),
  1066 => (x"fa",x"ff",x"fe",x"49"),
  1067 => (x"74",x"87",x"d8",x"87"),
  1068 => (x"c2",x"93",x"de",x"4b"),
  1069 => (x"cb",x"83",x"f4",x"da"),
  1070 => (x"51",x"c0",x"49",x"a3"),
  1071 => (x"6e",x"73",x"84",x"c1"),
  1072 => (x"fe",x"49",x"cb",x"4a"),
  1073 => (x"c4",x"87",x"e0",x"ff"),
  1074 => (x"80",x"c1",x"48",x"66"),
  1075 => (x"c7",x"58",x"a6",x"c8"),
  1076 => (x"c5",x"c0",x"03",x"ac"),
  1077 => (x"fc",x"05",x"6e",x"87"),
  1078 => (x"48",x"74",x"87",x"e4"),
  1079 => (x"e7",x"f5",x"8e",x"f4"),
  1080 => (x"1e",x"73",x"1e",x"87"),
  1081 => (x"cb",x"49",x"4b",x"71"),
  1082 => (x"f4",x"dd",x"c1",x"91"),
  1083 => (x"4a",x"a1",x"c8",x"81"),
  1084 => (x"48",x"e0",x"dd",x"c1"),
  1085 => (x"a1",x"c9",x"50",x"12"),
  1086 => (x"fb",x"f3",x"c0",x"4a"),
  1087 => (x"ca",x"50",x"12",x"48"),
  1088 => (x"e1",x"dd",x"c1",x"81"),
  1089 => (x"c1",x"50",x"11",x"48"),
  1090 => (x"bf",x"97",x"e1",x"dd"),
  1091 => (x"49",x"c0",x"1e",x"49"),
  1092 => (x"c2",x"87",x"fc",x"f5"),
  1093 => (x"de",x"48",x"c8",x"da"),
  1094 => (x"d5",x"49",x"c1",x"78"),
  1095 => (x"f4",x"26",x"87",x"ed"),
  1096 => (x"5e",x"0e",x"87",x"ea"),
  1097 => (x"0e",x"5d",x"5c",x"5b"),
  1098 => (x"4d",x"71",x"86",x"f4"),
  1099 => (x"c1",x"91",x"cb",x"49"),
  1100 => (x"c8",x"81",x"f4",x"dd"),
  1101 => (x"a1",x"ca",x"4a",x"a1"),
  1102 => (x"48",x"a6",x"c4",x"7e"),
  1103 => (x"bf",x"d0",x"de",x"c2"),
  1104 => (x"bf",x"97",x"6e",x"78"),
  1105 => (x"4c",x"66",x"c4",x"4b"),
  1106 => (x"48",x"12",x"2c",x"73"),
  1107 => (x"70",x"58",x"a6",x"cc"),
  1108 => (x"c9",x"84",x"c1",x"9c"),
  1109 => (x"49",x"69",x"97",x"81"),
  1110 => (x"c2",x"04",x"ac",x"b7"),
  1111 => (x"6e",x"4c",x"c0",x"87"),
  1112 => (x"c8",x"4a",x"bf",x"97"),
  1113 => (x"31",x"72",x"49",x"66"),
  1114 => (x"66",x"c4",x"b9",x"ff"),
  1115 => (x"72",x"48",x"74",x"99"),
  1116 => (x"48",x"4a",x"70",x"30"),
  1117 => (x"de",x"c2",x"b0",x"71"),
  1118 => (x"e4",x"c0",x"58",x"d4"),
  1119 => (x"49",x"c0",x"87",x"d7"),
  1120 => (x"75",x"87",x"c8",x"d4"),
  1121 => (x"cc",x"f6",x"c0",x"49"),
  1122 => (x"f2",x"8e",x"f4",x"87"),
  1123 => (x"73",x"1e",x"87",x"fa"),
  1124 => (x"49",x"4b",x"71",x"1e"),
  1125 => (x"73",x"87",x"cb",x"fe"),
  1126 => (x"87",x"c6",x"fe",x"49"),
  1127 => (x"1e",x"87",x"ed",x"f2"),
  1128 => (x"4b",x"71",x"1e",x"73"),
  1129 => (x"02",x"4a",x"a3",x"c6"),
  1130 => (x"8a",x"c1",x"87",x"db"),
  1131 => (x"8a",x"87",x"d6",x"02"),
  1132 => (x"87",x"da",x"c1",x"02"),
  1133 => (x"fc",x"c0",x"02",x"8a"),
  1134 => (x"c0",x"02",x"8a",x"87"),
  1135 => (x"02",x"8a",x"87",x"e1"),
  1136 => (x"db",x"c1",x"87",x"cb"),
  1137 => (x"f6",x"49",x"c7",x"87"),
  1138 => (x"de",x"c1",x"87",x"c7"),
  1139 => (x"e0",x"da",x"c2",x"87"),
  1140 => (x"cb",x"c1",x"02",x"bf"),
  1141 => (x"88",x"c1",x"48",x"87"),
  1142 => (x"58",x"e4",x"da",x"c2"),
  1143 => (x"c2",x"87",x"c1",x"c1"),
  1144 => (x"02",x"bf",x"e4",x"da"),
  1145 => (x"c2",x"87",x"f9",x"c0"),
  1146 => (x"48",x"bf",x"e0",x"da"),
  1147 => (x"da",x"c2",x"80",x"c1"),
  1148 => (x"eb",x"c0",x"58",x"e4"),
  1149 => (x"e0",x"da",x"c2",x"87"),
  1150 => (x"89",x"c6",x"49",x"bf"),
  1151 => (x"59",x"e4",x"da",x"c2"),
  1152 => (x"03",x"a9",x"b7",x"c0"),
  1153 => (x"da",x"c2",x"87",x"da"),
  1154 => (x"78",x"c0",x"48",x"e0"),
  1155 => (x"da",x"c2",x"87",x"d2"),
  1156 => (x"cb",x"02",x"bf",x"e4"),
  1157 => (x"e0",x"da",x"c2",x"87"),
  1158 => (x"80",x"c6",x"48",x"bf"),
  1159 => (x"58",x"e4",x"da",x"c2"),
  1160 => (x"e6",x"d1",x"49",x"c0"),
  1161 => (x"c0",x"49",x"73",x"87"),
  1162 => (x"f0",x"87",x"ea",x"f3"),
  1163 => (x"5e",x"0e",x"87",x"de"),
  1164 => (x"0e",x"5d",x"5c",x"5b"),
  1165 => (x"dc",x"86",x"d4",x"ff"),
  1166 => (x"a6",x"c8",x"59",x"a6"),
  1167 => (x"c4",x"78",x"c0",x"48"),
  1168 => (x"66",x"c0",x"c1",x"80"),
  1169 => (x"c1",x"80",x"c4",x"78"),
  1170 => (x"c1",x"80",x"c4",x"78"),
  1171 => (x"e4",x"da",x"c2",x"78"),
  1172 => (x"c2",x"78",x"c1",x"48"),
  1173 => (x"48",x"bf",x"c8",x"da"),
  1174 => (x"c9",x"05",x"a8",x"de"),
  1175 => (x"87",x"f8",x"f4",x"87"),
  1176 => (x"cf",x"58",x"a6",x"cc"),
  1177 => (x"e3",x"e4",x"87",x"e4"),
  1178 => (x"87",x"c5",x"e5",x"87"),
  1179 => (x"70",x"87",x"d2",x"e4"),
  1180 => (x"ac",x"fb",x"c0",x"4c"),
  1181 => (x"87",x"fb",x"c1",x"02"),
  1182 => (x"c1",x"05",x"66",x"d8"),
  1183 => (x"fc",x"c0",x"87",x"ed"),
  1184 => (x"82",x"c4",x"4a",x"66"),
  1185 => (x"1e",x"72",x"7e",x"6a"),
  1186 => (x"48",x"ff",x"d9",x"c1"),
  1187 => (x"c8",x"49",x"66",x"c4"),
  1188 => (x"41",x"20",x"4a",x"a1"),
  1189 => (x"f9",x"05",x"aa",x"71"),
  1190 => (x"26",x"51",x"10",x"87"),
  1191 => (x"66",x"fc",x"c0",x"4a"),
  1192 => (x"e1",x"c3",x"c1",x"48"),
  1193 => (x"c7",x"49",x"6a",x"78"),
  1194 => (x"c0",x"51",x"74",x"81"),
  1195 => (x"c8",x"49",x"66",x"fc"),
  1196 => (x"c0",x"51",x"c1",x"81"),
  1197 => (x"c9",x"49",x"66",x"fc"),
  1198 => (x"c0",x"51",x"c0",x"81"),
  1199 => (x"ca",x"49",x"66",x"fc"),
  1200 => (x"c1",x"51",x"c0",x"81"),
  1201 => (x"6a",x"1e",x"d8",x"1e"),
  1202 => (x"e3",x"81",x"c8",x"49"),
  1203 => (x"86",x"c8",x"87",x"f7"),
  1204 => (x"48",x"66",x"c0",x"c1"),
  1205 => (x"c7",x"01",x"a8",x"c0"),
  1206 => (x"48",x"a6",x"c8",x"87"),
  1207 => (x"87",x"ce",x"78",x"c1"),
  1208 => (x"48",x"66",x"c0",x"c1"),
  1209 => (x"a6",x"d0",x"88",x"c1"),
  1210 => (x"e3",x"87",x"c3",x"58"),
  1211 => (x"a6",x"d0",x"87",x"c3"),
  1212 => (x"74",x"78",x"c2",x"48"),
  1213 => (x"cd",x"cd",x"02",x"9c"),
  1214 => (x"48",x"66",x"c8",x"87"),
  1215 => (x"a8",x"66",x"c4",x"c1"),
  1216 => (x"87",x"c2",x"cd",x"03"),
  1217 => (x"c0",x"48",x"a6",x"dc"),
  1218 => (x"c0",x"80",x"e8",x"78"),
  1219 => (x"87",x"f1",x"e1",x"78"),
  1220 => (x"d0",x"c1",x"4c",x"70"),
  1221 => (x"d5",x"c2",x"05",x"ac"),
  1222 => (x"7e",x"66",x"c4",x"87"),
  1223 => (x"c8",x"87",x"d5",x"e4"),
  1224 => (x"dc",x"e1",x"58",x"a6"),
  1225 => (x"c0",x"4c",x"70",x"87"),
  1226 => (x"c1",x"05",x"ac",x"ec"),
  1227 => (x"66",x"c8",x"87",x"eb"),
  1228 => (x"c0",x"91",x"cb",x"49"),
  1229 => (x"c4",x"81",x"66",x"fc"),
  1230 => (x"4d",x"6a",x"4a",x"a1"),
  1231 => (x"c4",x"4a",x"a1",x"c8"),
  1232 => (x"fd",x"c0",x"52",x"66"),
  1233 => (x"f8",x"e0",x"79",x"d1"),
  1234 => (x"9c",x"4c",x"70",x"87"),
  1235 => (x"c0",x"87",x"d8",x"02"),
  1236 => (x"d2",x"02",x"ac",x"fb"),
  1237 => (x"e0",x"55",x"74",x"87"),
  1238 => (x"4c",x"70",x"87",x"e7"),
  1239 => (x"87",x"c7",x"02",x"9c"),
  1240 => (x"05",x"ac",x"fb",x"c0"),
  1241 => (x"c0",x"87",x"ee",x"ff"),
  1242 => (x"c1",x"c2",x"55",x"e0"),
  1243 => (x"7d",x"97",x"c0",x"55"),
  1244 => (x"6e",x"48",x"66",x"d8"),
  1245 => (x"87",x"db",x"05",x"a8"),
  1246 => (x"cc",x"48",x"66",x"c8"),
  1247 => (x"ca",x"04",x"a8",x"66"),
  1248 => (x"48",x"66",x"c8",x"87"),
  1249 => (x"a6",x"cc",x"80",x"c1"),
  1250 => (x"cc",x"87",x"c8",x"58"),
  1251 => (x"88",x"c1",x"48",x"66"),
  1252 => (x"ff",x"58",x"a6",x"d0"),
  1253 => (x"70",x"87",x"ea",x"df"),
  1254 => (x"ac",x"d0",x"c1",x"4c"),
  1255 => (x"d4",x"87",x"c8",x"05"),
  1256 => (x"80",x"c1",x"48",x"66"),
  1257 => (x"c1",x"58",x"a6",x"d8"),
  1258 => (x"fd",x"02",x"ac",x"d0"),
  1259 => (x"66",x"c4",x"87",x"eb"),
  1260 => (x"a8",x"66",x"d8",x"48"),
  1261 => (x"87",x"e0",x"c9",x"05"),
  1262 => (x"48",x"a6",x"e0",x"c0"),
  1263 => (x"48",x"74",x"78",x"c0"),
  1264 => (x"70",x"88",x"fb",x"c0"),
  1265 => (x"02",x"98",x"48",x"7e"),
  1266 => (x"48",x"87",x"e2",x"c9"),
  1267 => (x"7e",x"70",x"88",x"cb"),
  1268 => (x"c1",x"02",x"98",x"48"),
  1269 => (x"c9",x"48",x"87",x"cd"),
  1270 => (x"48",x"7e",x"70",x"88"),
  1271 => (x"fe",x"c3",x"02",x"98"),
  1272 => (x"88",x"c4",x"48",x"87"),
  1273 => (x"98",x"48",x"7e",x"70"),
  1274 => (x"48",x"87",x"ce",x"02"),
  1275 => (x"7e",x"70",x"88",x"c1"),
  1276 => (x"c3",x"02",x"98",x"48"),
  1277 => (x"d6",x"c8",x"87",x"e9"),
  1278 => (x"48",x"a6",x"dc",x"87"),
  1279 => (x"ff",x"78",x"f0",x"c0"),
  1280 => (x"70",x"87",x"fe",x"dd"),
  1281 => (x"ac",x"ec",x"c0",x"4c"),
  1282 => (x"87",x"c4",x"c0",x"02"),
  1283 => (x"5c",x"a6",x"e0",x"c0"),
  1284 => (x"02",x"ac",x"ec",x"c0"),
  1285 => (x"dd",x"ff",x"87",x"cd"),
  1286 => (x"4c",x"70",x"87",x"e7"),
  1287 => (x"05",x"ac",x"ec",x"c0"),
  1288 => (x"c0",x"87",x"f3",x"ff"),
  1289 => (x"c0",x"02",x"ac",x"ec"),
  1290 => (x"dd",x"ff",x"87",x"c4"),
  1291 => (x"1e",x"c0",x"87",x"d3"),
  1292 => (x"66",x"d0",x"1e",x"ca"),
  1293 => (x"c1",x"91",x"cb",x"49"),
  1294 => (x"71",x"48",x"66",x"c4"),
  1295 => (x"58",x"a6",x"cc",x"80"),
  1296 => (x"c4",x"48",x"66",x"c8"),
  1297 => (x"58",x"a6",x"d0",x"80"),
  1298 => (x"49",x"bf",x"66",x"cc"),
  1299 => (x"87",x"f5",x"dd",x"ff"),
  1300 => (x"1e",x"de",x"1e",x"c1"),
  1301 => (x"49",x"bf",x"66",x"d4"),
  1302 => (x"87",x"e9",x"dd",x"ff"),
  1303 => (x"49",x"70",x"86",x"d0"),
  1304 => (x"88",x"08",x"c0",x"48"),
  1305 => (x"58",x"a6",x"e8",x"c0"),
  1306 => (x"c0",x"06",x"a8",x"c0"),
  1307 => (x"e4",x"c0",x"87",x"ee"),
  1308 => (x"a8",x"dd",x"48",x"66"),
  1309 => (x"87",x"e4",x"c0",x"03"),
  1310 => (x"49",x"bf",x"66",x"c4"),
  1311 => (x"81",x"66",x"e4",x"c0"),
  1312 => (x"c0",x"51",x"e0",x"c0"),
  1313 => (x"c1",x"49",x"66",x"e4"),
  1314 => (x"bf",x"66",x"c4",x"81"),
  1315 => (x"51",x"c1",x"c2",x"81"),
  1316 => (x"49",x"66",x"e4",x"c0"),
  1317 => (x"66",x"c4",x"81",x"c2"),
  1318 => (x"51",x"c0",x"81",x"bf"),
  1319 => (x"c3",x"c1",x"48",x"6e"),
  1320 => (x"49",x"6e",x"78",x"e1"),
  1321 => (x"66",x"d0",x"81",x"c8"),
  1322 => (x"c9",x"49",x"6e",x"51"),
  1323 => (x"51",x"66",x"d4",x"81"),
  1324 => (x"81",x"ca",x"49",x"6e"),
  1325 => (x"d0",x"51",x"66",x"dc"),
  1326 => (x"80",x"c1",x"48",x"66"),
  1327 => (x"c8",x"58",x"a6",x"d4"),
  1328 => (x"66",x"cc",x"48",x"66"),
  1329 => (x"cb",x"c0",x"04",x"a8"),
  1330 => (x"48",x"66",x"c8",x"87"),
  1331 => (x"a6",x"cc",x"80",x"c1"),
  1332 => (x"87",x"d9",x"c5",x"58"),
  1333 => (x"c1",x"48",x"66",x"cc"),
  1334 => (x"58",x"a6",x"d0",x"88"),
  1335 => (x"ff",x"87",x"ce",x"c5"),
  1336 => (x"c0",x"87",x"d1",x"dd"),
  1337 => (x"ff",x"58",x"a6",x"e8"),
  1338 => (x"c0",x"87",x"c9",x"dd"),
  1339 => (x"c0",x"58",x"a6",x"e0"),
  1340 => (x"c0",x"05",x"a8",x"ec"),
  1341 => (x"a6",x"dc",x"87",x"ca"),
  1342 => (x"66",x"e4",x"c0",x"48"),
  1343 => (x"87",x"c4",x"c0",x"78"),
  1344 => (x"87",x"fd",x"d9",x"ff"),
  1345 => (x"cb",x"49",x"66",x"c8"),
  1346 => (x"66",x"fc",x"c0",x"91"),
  1347 => (x"70",x"80",x"71",x"48"),
  1348 => (x"82",x"c8",x"4a",x"7e"),
  1349 => (x"81",x"ca",x"49",x"6e"),
  1350 => (x"51",x"66",x"e4",x"c0"),
  1351 => (x"c1",x"49",x"66",x"dc"),
  1352 => (x"66",x"e4",x"c0",x"81"),
  1353 => (x"71",x"48",x"c1",x"89"),
  1354 => (x"c1",x"49",x"70",x"30"),
  1355 => (x"7a",x"97",x"71",x"89"),
  1356 => (x"bf",x"d0",x"de",x"c2"),
  1357 => (x"66",x"e4",x"c0",x"49"),
  1358 => (x"4a",x"6a",x"97",x"29"),
  1359 => (x"c0",x"98",x"71",x"48"),
  1360 => (x"6e",x"58",x"a6",x"ec"),
  1361 => (x"69",x"81",x"c4",x"49"),
  1362 => (x"48",x"66",x"d8",x"4d"),
  1363 => (x"02",x"a8",x"66",x"c4"),
  1364 => (x"c4",x"87",x"c8",x"c0"),
  1365 => (x"78",x"c0",x"48",x"a6"),
  1366 => (x"c4",x"87",x"c5",x"c0"),
  1367 => (x"78",x"c1",x"48",x"a6"),
  1368 => (x"c0",x"1e",x"66",x"c4"),
  1369 => (x"49",x"75",x"1e",x"e0"),
  1370 => (x"87",x"d9",x"d9",x"ff"),
  1371 => (x"4c",x"70",x"86",x"c8"),
  1372 => (x"06",x"ac",x"b7",x"c0"),
  1373 => (x"74",x"87",x"d4",x"c1"),
  1374 => (x"49",x"e0",x"c0",x"85"),
  1375 => (x"4b",x"75",x"89",x"74"),
  1376 => (x"4a",x"c8",x"da",x"c1"),
  1377 => (x"de",x"ec",x"fe",x"71"),
  1378 => (x"c0",x"85",x"c2",x"87"),
  1379 => (x"c1",x"48",x"66",x"e0"),
  1380 => (x"a6",x"e4",x"c0",x"80"),
  1381 => (x"66",x"e8",x"c0",x"58"),
  1382 => (x"70",x"81",x"c1",x"49"),
  1383 => (x"c8",x"c0",x"02",x"a9"),
  1384 => (x"48",x"a6",x"c4",x"87"),
  1385 => (x"c5",x"c0",x"78",x"c0"),
  1386 => (x"48",x"a6",x"c4",x"87"),
  1387 => (x"66",x"c4",x"78",x"c1"),
  1388 => (x"49",x"a4",x"c2",x"1e"),
  1389 => (x"71",x"48",x"e0",x"c0"),
  1390 => (x"1e",x"49",x"70",x"88"),
  1391 => (x"d8",x"ff",x"49",x"75"),
  1392 => (x"86",x"c8",x"87",x"c3"),
  1393 => (x"01",x"a8",x"b7",x"c0"),
  1394 => (x"c0",x"87",x"c0",x"ff"),
  1395 => (x"c0",x"02",x"66",x"e0"),
  1396 => (x"49",x"6e",x"87",x"d1"),
  1397 => (x"e0",x"c0",x"81",x"c9"),
  1398 => (x"48",x"6e",x"51",x"66"),
  1399 => (x"78",x"e2",x"c4",x"c1"),
  1400 => (x"6e",x"87",x"cc",x"c0"),
  1401 => (x"c2",x"81",x"c9",x"49"),
  1402 => (x"c1",x"48",x"6e",x"51"),
  1403 => (x"c8",x"78",x"ce",x"c6"),
  1404 => (x"66",x"cc",x"48",x"66"),
  1405 => (x"cb",x"c0",x"04",x"a8"),
  1406 => (x"48",x"66",x"c8",x"87"),
  1407 => (x"a6",x"cc",x"80",x"c1"),
  1408 => (x"87",x"e9",x"c0",x"58"),
  1409 => (x"c1",x"48",x"66",x"cc"),
  1410 => (x"58",x"a6",x"d0",x"88"),
  1411 => (x"ff",x"87",x"de",x"c0"),
  1412 => (x"70",x"87",x"de",x"d6"),
  1413 => (x"87",x"d5",x"c0",x"4c"),
  1414 => (x"05",x"ac",x"c6",x"c1"),
  1415 => (x"d0",x"87",x"c8",x"c0"),
  1416 => (x"80",x"c1",x"48",x"66"),
  1417 => (x"ff",x"58",x"a6",x"d4"),
  1418 => (x"70",x"87",x"c6",x"d6"),
  1419 => (x"48",x"66",x"d4",x"4c"),
  1420 => (x"a6",x"d8",x"80",x"c1"),
  1421 => (x"02",x"9c",x"74",x"58"),
  1422 => (x"c8",x"87",x"cb",x"c0"),
  1423 => (x"c4",x"c1",x"48",x"66"),
  1424 => (x"f2",x"04",x"a8",x"66"),
  1425 => (x"d5",x"ff",x"87",x"fe"),
  1426 => (x"66",x"c8",x"87",x"de"),
  1427 => (x"03",x"a8",x"c7",x"48"),
  1428 => (x"c2",x"87",x"e5",x"c0"),
  1429 => (x"c0",x"48",x"e4",x"da"),
  1430 => (x"49",x"66",x"c8",x"78"),
  1431 => (x"fc",x"c0",x"91",x"cb"),
  1432 => (x"a1",x"c4",x"81",x"66"),
  1433 => (x"c0",x"4a",x"6a",x"4a"),
  1434 => (x"66",x"c8",x"79",x"52"),
  1435 => (x"cc",x"80",x"c1",x"48"),
  1436 => (x"a8",x"c7",x"58",x"a6"),
  1437 => (x"87",x"db",x"ff",x"04"),
  1438 => (x"ff",x"8e",x"d4",x"ff"),
  1439 => (x"4c",x"87",x"c9",x"df"),
  1440 => (x"20",x"64",x"61",x"6f"),
  1441 => (x"00",x"20",x"2e",x"2a"),
  1442 => (x"1e",x"00",x"20",x"3a"),
  1443 => (x"4b",x"71",x"1e",x"73"),
  1444 => (x"87",x"c6",x"02",x"9b"),
  1445 => (x"48",x"e0",x"da",x"c2"),
  1446 => (x"1e",x"c7",x"78",x"c0"),
  1447 => (x"bf",x"e0",x"da",x"c2"),
  1448 => (x"f4",x"dd",x"c1",x"1e"),
  1449 => (x"c8",x"da",x"c2",x"1e"),
  1450 => (x"c1",x"ee",x"49",x"bf"),
  1451 => (x"c2",x"86",x"cc",x"87"),
  1452 => (x"49",x"bf",x"c8",x"da"),
  1453 => (x"73",x"87",x"f9",x"e2"),
  1454 => (x"87",x"c8",x"02",x"9b"),
  1455 => (x"49",x"f4",x"dd",x"c1"),
  1456 => (x"87",x"e3",x"e2",x"c0"),
  1457 => (x"87",x"c4",x"de",x"ff"),
  1458 => (x"e0",x"dd",x"c1",x"1e"),
  1459 => (x"c1",x"50",x"c0",x"48"),
  1460 => (x"49",x"bf",x"d7",x"df"),
  1461 => (x"87",x"e4",x"d8",x"ff"),
  1462 => (x"4f",x"26",x"48",x"c0"),
  1463 => (x"87",x"de",x"c7",x"1e"),
  1464 => (x"e6",x"fe",x"49",x"c1"),
  1465 => (x"c7",x"ef",x"fe",x"87"),
  1466 => (x"02",x"98",x"70",x"87"),
  1467 => (x"f6",x"fe",x"87",x"cd"),
  1468 => (x"98",x"70",x"87",x"e1"),
  1469 => (x"c1",x"87",x"c4",x"02"),
  1470 => (x"c0",x"87",x"c2",x"4a"),
  1471 => (x"05",x"9a",x"72",x"4a"),
  1472 => (x"1e",x"c0",x"87",x"ce"),
  1473 => (x"49",x"f7",x"dc",x"c1"),
  1474 => (x"87",x"de",x"ee",x"c0"),
  1475 => (x"87",x"fe",x"86",x"c4"),
  1476 => (x"48",x"e0",x"da",x"c2"),
  1477 => (x"da",x"c2",x"78",x"c0"),
  1478 => (x"78",x"c0",x"48",x"c8"),
  1479 => (x"c2",x"dd",x"c1",x"1e"),
  1480 => (x"c5",x"ee",x"c0",x"49"),
  1481 => (x"fe",x"1e",x"c0",x"87"),
  1482 => (x"49",x"70",x"87",x"de"),
  1483 => (x"87",x"fa",x"ed",x"c0"),
  1484 => (x"f8",x"87",x"ca",x"c3"),
  1485 => (x"53",x"4f",x"26",x"8e"),
  1486 => (x"61",x"66",x"20",x"44"),
  1487 => (x"64",x"65",x"6c",x"69"),
  1488 => (x"6f",x"42",x"00",x"2e"),
  1489 => (x"6e",x"69",x"74",x"6f"),
  1490 => (x"2e",x"2e",x"2e",x"67"),
  1491 => (x"e2",x"c0",x"1e",x"00"),
  1492 => (x"87",x"fa",x"87",x"d2"),
  1493 => (x"fe",x"1e",x"4f",x"26"),
  1494 => (x"87",x"f1",x"87",x"c2"),
  1495 => (x"4f",x"26",x"48",x"c0"),
  1496 => (x"00",x"01",x"00",x"00"),
  1497 => (x"20",x"80",x"00",x"00"),
  1498 => (x"74",x"69",x"78",x"45"),
  1499 => (x"42",x"20",x"80",x"00"),
  1500 => (x"00",x"6b",x"63",x"61"),
  1501 => (x"00",x"00",x"0e",x"9e"),
  1502 => (x"00",x"00",x"26",x"b4"),
  1503 => (x"9e",x"00",x"00",x"00"),
  1504 => (x"d2",x"00",x"00",x"0e"),
  1505 => (x"00",x"00",x"00",x"26"),
  1506 => (x"0e",x"9e",x"00",x"00"),
  1507 => (x"26",x"f0",x"00",x"00"),
  1508 => (x"00",x"00",x"00",x"00"),
  1509 => (x"00",x"0e",x"9e",x"00"),
  1510 => (x"00",x"27",x"0e",x"00"),
  1511 => (x"00",x"00",x"00",x"00"),
  1512 => (x"00",x"00",x"0e",x"9e"),
  1513 => (x"00",x"00",x"27",x"2c"),
  1514 => (x"9e",x"00",x"00",x"00"),
  1515 => (x"4a",x"00",x"00",x"0e"),
  1516 => (x"00",x"00",x"00",x"27"),
  1517 => (x"0e",x"9e",x"00",x"00"),
  1518 => (x"27",x"68",x"00",x"00"),
  1519 => (x"00",x"00",x"00",x"00"),
  1520 => (x"00",x"0f",x"51",x"00"),
  1521 => (x"00",x"00",x"00",x"00"),
  1522 => (x"00",x"00",x"00",x"00"),
  1523 => (x"00",x"00",x"11",x"9f"),
  1524 => (x"00",x"00",x"00",x"00"),
  1525 => (x"db",x"00",x"00",x"00"),
  1526 => (x"42",x"00",x"00",x"17"),
  1527 => (x"20",x"54",x"4f",x"4f"),
  1528 => (x"52",x"20",x"20",x"20"),
  1529 => (x"1e",x"00",x"4d",x"4f"),
  1530 => (x"c0",x"48",x"f0",x"fe"),
  1531 => (x"79",x"09",x"cd",x"78"),
  1532 => (x"1e",x"4f",x"26",x"09"),
  1533 => (x"bf",x"f0",x"fe",x"1e"),
  1534 => (x"26",x"26",x"48",x"7e"),
  1535 => (x"f0",x"fe",x"1e",x"4f"),
  1536 => (x"26",x"78",x"c1",x"48"),
  1537 => (x"f0",x"fe",x"1e",x"4f"),
  1538 => (x"26",x"78",x"c0",x"48"),
  1539 => (x"4a",x"71",x"1e",x"4f"),
  1540 => (x"26",x"52",x"52",x"c0"),
  1541 => (x"5b",x"5e",x"0e",x"4f"),
  1542 => (x"f4",x"0e",x"5d",x"5c"),
  1543 => (x"97",x"4d",x"71",x"86"),
  1544 => (x"a5",x"c1",x"7e",x"6d"),
  1545 => (x"48",x"6c",x"97",x"4c"),
  1546 => (x"6e",x"58",x"a6",x"c8"),
  1547 => (x"a8",x"66",x"c4",x"48"),
  1548 => (x"ff",x"87",x"c5",x"05"),
  1549 => (x"87",x"e6",x"c0",x"48"),
  1550 => (x"c2",x"87",x"ca",x"ff"),
  1551 => (x"6c",x"97",x"49",x"a5"),
  1552 => (x"4b",x"a3",x"71",x"4b"),
  1553 => (x"97",x"4b",x"6b",x"97"),
  1554 => (x"48",x"6e",x"7e",x"6c"),
  1555 => (x"a6",x"c8",x"80",x"c1"),
  1556 => (x"cc",x"98",x"c7",x"58"),
  1557 => (x"97",x"70",x"58",x"a6"),
  1558 => (x"87",x"e1",x"fe",x"7c"),
  1559 => (x"8e",x"f4",x"48",x"73"),
  1560 => (x"4c",x"26",x"4d",x"26"),
  1561 => (x"4f",x"26",x"4b",x"26"),
  1562 => (x"5c",x"5b",x"5e",x"0e"),
  1563 => (x"71",x"86",x"f4",x"0e"),
  1564 => (x"4a",x"66",x"d8",x"4c"),
  1565 => (x"c2",x"9a",x"ff",x"c3"),
  1566 => (x"6c",x"97",x"4b",x"a4"),
  1567 => (x"49",x"a1",x"73",x"49"),
  1568 => (x"6c",x"97",x"51",x"72"),
  1569 => (x"c1",x"48",x"6e",x"7e"),
  1570 => (x"58",x"a6",x"c8",x"80"),
  1571 => (x"a6",x"cc",x"98",x"c7"),
  1572 => (x"f4",x"54",x"70",x"58"),
  1573 => (x"87",x"ca",x"ff",x"8e"),
  1574 => (x"e8",x"fd",x"1e",x"1e"),
  1575 => (x"4a",x"bf",x"e0",x"87"),
  1576 => (x"c0",x"e0",x"c0",x"49"),
  1577 => (x"87",x"cb",x"02",x"99"),
  1578 => (x"de",x"c2",x"1e",x"72"),
  1579 => (x"f7",x"fe",x"49",x"c6"),
  1580 => (x"fc",x"86",x"c4",x"87"),
  1581 => (x"7e",x"70",x"87",x"fd"),
  1582 => (x"26",x"87",x"c2",x"fd"),
  1583 => (x"c2",x"1e",x"4f",x"26"),
  1584 => (x"fd",x"49",x"c6",x"de"),
  1585 => (x"e2",x"c1",x"87",x"c7"),
  1586 => (x"da",x"fc",x"49",x"d8"),
  1587 => (x"87",x"ee",x"c3",x"87"),
  1588 => (x"5e",x"0e",x"4f",x"26"),
  1589 => (x"0e",x"5d",x"5c",x"5b"),
  1590 => (x"de",x"c2",x"4d",x"71"),
  1591 => (x"f4",x"fc",x"49",x"c6"),
  1592 => (x"c0",x"4b",x"70",x"87"),
  1593 => (x"c3",x"04",x"ab",x"b7"),
  1594 => (x"f0",x"c3",x"87",x"c2"),
  1595 => (x"87",x"c9",x"05",x"ab"),
  1596 => (x"48",x"f6",x"e6",x"c1"),
  1597 => (x"e3",x"c2",x"78",x"c1"),
  1598 => (x"ab",x"e0",x"c3",x"87"),
  1599 => (x"c1",x"87",x"c9",x"05"),
  1600 => (x"c1",x"48",x"fa",x"e6"),
  1601 => (x"87",x"d4",x"c2",x"78"),
  1602 => (x"bf",x"fa",x"e6",x"c1"),
  1603 => (x"c2",x"87",x"c6",x"02"),
  1604 => (x"c2",x"4c",x"a3",x"c0"),
  1605 => (x"c1",x"4c",x"73",x"87"),
  1606 => (x"02",x"bf",x"f6",x"e6"),
  1607 => (x"74",x"87",x"e0",x"c0"),
  1608 => (x"29",x"b7",x"c4",x"49"),
  1609 => (x"cd",x"e8",x"c1",x"91"),
  1610 => (x"cf",x"4a",x"74",x"81"),
  1611 => (x"c1",x"92",x"c2",x"9a"),
  1612 => (x"70",x"30",x"72",x"48"),
  1613 => (x"72",x"ba",x"ff",x"4a"),
  1614 => (x"70",x"98",x"69",x"48"),
  1615 => (x"74",x"87",x"db",x"79"),
  1616 => (x"29",x"b7",x"c4",x"49"),
  1617 => (x"cd",x"e8",x"c1",x"91"),
  1618 => (x"cf",x"4a",x"74",x"81"),
  1619 => (x"c3",x"92",x"c2",x"9a"),
  1620 => (x"70",x"30",x"72",x"48"),
  1621 => (x"b0",x"69",x"48",x"4a"),
  1622 => (x"9d",x"75",x"79",x"70"),
  1623 => (x"87",x"f0",x"c0",x"05"),
  1624 => (x"c8",x"48",x"d0",x"ff"),
  1625 => (x"d4",x"ff",x"78",x"e1"),
  1626 => (x"c1",x"78",x"c5",x"48"),
  1627 => (x"02",x"bf",x"fa",x"e6"),
  1628 => (x"e0",x"c3",x"87",x"c3"),
  1629 => (x"f6",x"e6",x"c1",x"78"),
  1630 => (x"87",x"c6",x"02",x"bf"),
  1631 => (x"c3",x"48",x"d4",x"ff"),
  1632 => (x"d4",x"ff",x"78",x"f0"),
  1633 => (x"ff",x"0b",x"7b",x"0b"),
  1634 => (x"e1",x"c8",x"48",x"d0"),
  1635 => (x"78",x"e0",x"c0",x"78"),
  1636 => (x"48",x"fa",x"e6",x"c1"),
  1637 => (x"e6",x"c1",x"78",x"c0"),
  1638 => (x"78",x"c0",x"48",x"f6"),
  1639 => (x"49",x"c6",x"de",x"c2"),
  1640 => (x"70",x"87",x"f2",x"f9"),
  1641 => (x"ab",x"b7",x"c0",x"4b"),
  1642 => (x"87",x"fe",x"fc",x"03"),
  1643 => (x"4d",x"26",x"48",x"c0"),
  1644 => (x"4b",x"26",x"4c",x"26"),
  1645 => (x"00",x"00",x"4f",x"26"),
  1646 => (x"00",x"00",x"00",x"00"),
  1647 => (x"c0",x"1e",x"00",x"00"),
  1648 => (x"c4",x"49",x"72",x"4a"),
  1649 => (x"cd",x"e8",x"c1",x"91"),
  1650 => (x"c1",x"79",x"c0",x"81"),
  1651 => (x"aa",x"b7",x"d0",x"82"),
  1652 => (x"26",x"87",x"ee",x"04"),
  1653 => (x"5b",x"5e",x"0e",x"4f"),
  1654 => (x"71",x"0e",x"5d",x"5c"),
  1655 => (x"87",x"e5",x"f8",x"4d"),
  1656 => (x"b7",x"c4",x"4a",x"75"),
  1657 => (x"e8",x"c1",x"92",x"2a"),
  1658 => (x"4c",x"75",x"82",x"cd"),
  1659 => (x"94",x"c2",x"9c",x"cf"),
  1660 => (x"74",x"4b",x"49",x"6a"),
  1661 => (x"c2",x"9b",x"c3",x"2b"),
  1662 => (x"70",x"30",x"74",x"48"),
  1663 => (x"74",x"bc",x"ff",x"4c"),
  1664 => (x"70",x"98",x"71",x"48"),
  1665 => (x"87",x"f5",x"f7",x"7a"),
  1666 => (x"e1",x"fe",x"48",x"73"),
  1667 => (x"00",x"00",x"00",x"87"),
  1668 => (x"00",x"00",x"00",x"00"),
  1669 => (x"00",x"00",x"00",x"00"),
  1670 => (x"00",x"00",x"00",x"00"),
  1671 => (x"00",x"00",x"00",x"00"),
  1672 => (x"00",x"00",x"00",x"00"),
  1673 => (x"00",x"00",x"00",x"00"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"00",x"00",x"00",x"00"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"00",x"00",x"00",x"00"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"00",x"00",x"00"),
  1682 => (x"00",x"00",x"00",x"00"),
  1683 => (x"d0",x"ff",x"1e",x"00"),
  1684 => (x"78",x"e1",x"c8",x"48"),
  1685 => (x"d4",x"ff",x"48",x"71"),
  1686 => (x"66",x"c4",x"78",x"08"),
  1687 => (x"08",x"d4",x"ff",x"48"),
  1688 => (x"1e",x"4f",x"26",x"78"),
  1689 => (x"66",x"c4",x"4a",x"71"),
  1690 => (x"49",x"72",x"1e",x"49"),
  1691 => (x"ff",x"87",x"de",x"ff"),
  1692 => (x"e0",x"c0",x"48",x"d0"),
  1693 => (x"4f",x"26",x"26",x"78"),
  1694 => (x"71",x"1e",x"73",x"1e"),
  1695 => (x"49",x"66",x"c8",x"4b"),
  1696 => (x"c1",x"4a",x"73",x"1e"),
  1697 => (x"ff",x"49",x"a2",x"e0"),
  1698 => (x"c4",x"26",x"87",x"d9"),
  1699 => (x"26",x"4d",x"26",x"87"),
  1700 => (x"26",x"4b",x"26",x"4c"),
  1701 => (x"d4",x"ff",x"1e",x"4f"),
  1702 => (x"7a",x"ff",x"c3",x"4a"),
  1703 => (x"c0",x"48",x"d0",x"ff"),
  1704 => (x"7a",x"de",x"78",x"e1"),
  1705 => (x"bf",x"d0",x"de",x"c2"),
  1706 => (x"c8",x"48",x"49",x"7a"),
  1707 => (x"71",x"7a",x"70",x"28"),
  1708 => (x"70",x"28",x"d0",x"48"),
  1709 => (x"d8",x"48",x"71",x"7a"),
  1710 => (x"ff",x"7a",x"70",x"28"),
  1711 => (x"e0",x"c0",x"48",x"d0"),
  1712 => (x"1e",x"4f",x"26",x"78"),
  1713 => (x"c8",x"48",x"d0",x"ff"),
  1714 => (x"48",x"71",x"78",x"c9"),
  1715 => (x"78",x"08",x"d4",x"ff"),
  1716 => (x"71",x"1e",x"4f",x"26"),
  1717 => (x"87",x"eb",x"49",x"4a"),
  1718 => (x"c8",x"48",x"d0",x"ff"),
  1719 => (x"1e",x"4f",x"26",x"78"),
  1720 => (x"4b",x"71",x"1e",x"73"),
  1721 => (x"bf",x"e0",x"de",x"c2"),
  1722 => (x"c2",x"87",x"c3",x"02"),
  1723 => (x"d0",x"ff",x"87",x"eb"),
  1724 => (x"78",x"c9",x"c8",x"48"),
  1725 => (x"e0",x"c0",x"48",x"73"),
  1726 => (x"08",x"d4",x"ff",x"b0"),
  1727 => (x"d4",x"de",x"c2",x"78"),
  1728 => (x"c8",x"78",x"c0",x"48"),
  1729 => (x"87",x"c5",x"02",x"66"),
  1730 => (x"c2",x"49",x"ff",x"c3"),
  1731 => (x"c2",x"49",x"c0",x"87"),
  1732 => (x"cc",x"59",x"dc",x"de"),
  1733 => (x"87",x"c6",x"02",x"66"),
  1734 => (x"4a",x"d5",x"d5",x"c5"),
  1735 => (x"ff",x"cf",x"87",x"c4"),
  1736 => (x"de",x"c2",x"4a",x"ff"),
  1737 => (x"de",x"c2",x"5a",x"e0"),
  1738 => (x"78",x"c1",x"48",x"e0"),
  1739 => (x"4d",x"26",x"87",x"c4"),
  1740 => (x"4b",x"26",x"4c",x"26"),
  1741 => (x"5e",x"0e",x"4f",x"26"),
  1742 => (x"0e",x"5d",x"5c",x"5b"),
  1743 => (x"de",x"c2",x"4a",x"71"),
  1744 => (x"72",x"4c",x"bf",x"dc"),
  1745 => (x"87",x"cb",x"02",x"9a"),
  1746 => (x"c1",x"91",x"c8",x"49"),
  1747 => (x"71",x"4b",x"d5",x"eb"),
  1748 => (x"c1",x"87",x"c4",x"83"),
  1749 => (x"c0",x"4b",x"d5",x"ef"),
  1750 => (x"74",x"49",x"13",x"4d"),
  1751 => (x"d8",x"de",x"c2",x"99"),
  1752 => (x"b8",x"71",x"48",x"bf"),
  1753 => (x"78",x"08",x"d4",x"ff"),
  1754 => (x"85",x"2c",x"b7",x"c1"),
  1755 => (x"04",x"ad",x"b7",x"c8"),
  1756 => (x"de",x"c2",x"87",x"e7"),
  1757 => (x"c8",x"48",x"bf",x"d4"),
  1758 => (x"d8",x"de",x"c2",x"80"),
  1759 => (x"87",x"ee",x"fe",x"58"),
  1760 => (x"71",x"1e",x"73",x"1e"),
  1761 => (x"9a",x"4a",x"13",x"4b"),
  1762 => (x"72",x"87",x"cb",x"02"),
  1763 => (x"87",x"e6",x"fe",x"49"),
  1764 => (x"05",x"9a",x"4a",x"13"),
  1765 => (x"d9",x"fe",x"87",x"f5"),
  1766 => (x"de",x"c2",x"1e",x"87"),
  1767 => (x"c2",x"49",x"bf",x"d4"),
  1768 => (x"c1",x"48",x"d4",x"de"),
  1769 => (x"c0",x"c4",x"78",x"a1"),
  1770 => (x"db",x"03",x"a9",x"b7"),
  1771 => (x"48",x"d4",x"ff",x"87"),
  1772 => (x"bf",x"d8",x"de",x"c2"),
  1773 => (x"d4",x"de",x"c2",x"78"),
  1774 => (x"de",x"c2",x"49",x"bf"),
  1775 => (x"a1",x"c1",x"48",x"d4"),
  1776 => (x"b7",x"c0",x"c4",x"78"),
  1777 => (x"87",x"e5",x"04",x"a9"),
  1778 => (x"c8",x"48",x"d0",x"ff"),
  1779 => (x"e0",x"de",x"c2",x"78"),
  1780 => (x"26",x"78",x"c0",x"48"),
  1781 => (x"00",x"00",x"00",x"4f"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"5f",x"5f"),
  1785 => (x"03",x"03",x"00",x"00"),
  1786 => (x"00",x"03",x"03",x"00"),
  1787 => (x"7f",x"7f",x"14",x"00"),
  1788 => (x"14",x"7f",x"7f",x"14"),
  1789 => (x"2e",x"24",x"00",x"00"),
  1790 => (x"12",x"3a",x"6b",x"6b"),
  1791 => (x"36",x"6a",x"4c",x"00"),
  1792 => (x"32",x"56",x"6c",x"18"),
  1793 => (x"4f",x"7e",x"30",x"00"),
  1794 => (x"68",x"3a",x"77",x"59"),
  1795 => (x"04",x"00",x"00",x"40"),
  1796 => (x"00",x"00",x"03",x"07"),
  1797 => (x"1c",x"00",x"00",x"00"),
  1798 => (x"00",x"41",x"63",x"3e"),
  1799 => (x"41",x"00",x"00",x"00"),
  1800 => (x"00",x"1c",x"3e",x"63"),
  1801 => (x"3e",x"2a",x"08",x"00"),
  1802 => (x"2a",x"3e",x"1c",x"1c"),
  1803 => (x"08",x"08",x"00",x"08"),
  1804 => (x"08",x"08",x"3e",x"3e"),
  1805 => (x"80",x"00",x"00",x"00"),
  1806 => (x"00",x"00",x"60",x"e0"),
  1807 => (x"08",x"08",x"00",x"00"),
  1808 => (x"08",x"08",x"08",x"08"),
  1809 => (x"00",x"00",x"00",x"00"),
  1810 => (x"00",x"00",x"60",x"60"),
  1811 => (x"30",x"60",x"40",x"00"),
  1812 => (x"03",x"06",x"0c",x"18"),
  1813 => (x"7f",x"3e",x"00",x"01"),
  1814 => (x"3e",x"7f",x"4d",x"59"),
  1815 => (x"06",x"04",x"00",x"00"),
  1816 => (x"00",x"00",x"7f",x"7f"),
  1817 => (x"63",x"42",x"00",x"00"),
  1818 => (x"46",x"4f",x"59",x"71"),
  1819 => (x"63",x"22",x"00",x"00"),
  1820 => (x"36",x"7f",x"49",x"49"),
  1821 => (x"16",x"1c",x"18",x"00"),
  1822 => (x"10",x"7f",x"7f",x"13"),
  1823 => (x"67",x"27",x"00",x"00"),
  1824 => (x"39",x"7d",x"45",x"45"),
  1825 => (x"7e",x"3c",x"00",x"00"),
  1826 => (x"30",x"79",x"49",x"4b"),
  1827 => (x"01",x"01",x"00",x"00"),
  1828 => (x"07",x"0f",x"79",x"71"),
  1829 => (x"7f",x"36",x"00",x"00"),
  1830 => (x"36",x"7f",x"49",x"49"),
  1831 => (x"4f",x"06",x"00",x"00"),
  1832 => (x"1e",x"3f",x"69",x"49"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"00",x"00",x"66",x"66"),
  1835 => (x"80",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"66",x"e6"),
  1837 => (x"08",x"08",x"00",x"00"),
  1838 => (x"22",x"22",x"14",x"14"),
  1839 => (x"14",x"14",x"00",x"00"),
  1840 => (x"14",x"14",x"14",x"14"),
  1841 => (x"22",x"22",x"00",x"00"),
  1842 => (x"08",x"08",x"14",x"14"),
  1843 => (x"03",x"02",x"00",x"00"),
  1844 => (x"06",x"0f",x"59",x"51"),
  1845 => (x"41",x"7f",x"3e",x"00"),
  1846 => (x"1e",x"1f",x"55",x"5d"),
  1847 => (x"7f",x"7e",x"00",x"00"),
  1848 => (x"7e",x"7f",x"09",x"09"),
  1849 => (x"7f",x"7f",x"00",x"00"),
  1850 => (x"36",x"7f",x"49",x"49"),
  1851 => (x"3e",x"1c",x"00",x"00"),
  1852 => (x"41",x"41",x"41",x"63"),
  1853 => (x"7f",x"7f",x"00",x"00"),
  1854 => (x"1c",x"3e",x"63",x"41"),
  1855 => (x"7f",x"7f",x"00",x"00"),
  1856 => (x"41",x"41",x"49",x"49"),
  1857 => (x"7f",x"7f",x"00",x"00"),
  1858 => (x"01",x"01",x"09",x"09"),
  1859 => (x"7f",x"3e",x"00",x"00"),
  1860 => (x"7a",x"7b",x"49",x"41"),
  1861 => (x"7f",x"7f",x"00",x"00"),
  1862 => (x"7f",x"7f",x"08",x"08"),
  1863 => (x"41",x"00",x"00",x"00"),
  1864 => (x"00",x"41",x"7f",x"7f"),
  1865 => (x"60",x"20",x"00",x"00"),
  1866 => (x"3f",x"7f",x"40",x"40"),
  1867 => (x"08",x"7f",x"7f",x"00"),
  1868 => (x"41",x"63",x"36",x"1c"),
  1869 => (x"7f",x"7f",x"00",x"00"),
  1870 => (x"40",x"40",x"40",x"40"),
  1871 => (x"06",x"7f",x"7f",x"00"),
  1872 => (x"7f",x"7f",x"06",x"0c"),
  1873 => (x"06",x"7f",x"7f",x"00"),
  1874 => (x"7f",x"7f",x"18",x"0c"),
  1875 => (x"7f",x"3e",x"00",x"00"),
  1876 => (x"3e",x"7f",x"41",x"41"),
  1877 => (x"7f",x"7f",x"00",x"00"),
  1878 => (x"06",x"0f",x"09",x"09"),
  1879 => (x"41",x"7f",x"3e",x"00"),
  1880 => (x"40",x"7e",x"7f",x"61"),
  1881 => (x"7f",x"7f",x"00",x"00"),
  1882 => (x"66",x"7f",x"19",x"09"),
  1883 => (x"6f",x"26",x"00",x"00"),
  1884 => (x"32",x"7b",x"59",x"4d"),
  1885 => (x"01",x"01",x"00",x"00"),
  1886 => (x"01",x"01",x"7f",x"7f"),
  1887 => (x"7f",x"3f",x"00",x"00"),
  1888 => (x"3f",x"7f",x"40",x"40"),
  1889 => (x"3f",x"0f",x"00",x"00"),
  1890 => (x"0f",x"3f",x"70",x"70"),
  1891 => (x"30",x"7f",x"7f",x"00"),
  1892 => (x"7f",x"7f",x"30",x"18"),
  1893 => (x"36",x"63",x"41",x"00"),
  1894 => (x"63",x"36",x"1c",x"1c"),
  1895 => (x"06",x"03",x"01",x"41"),
  1896 => (x"03",x"06",x"7c",x"7c"),
  1897 => (x"59",x"71",x"61",x"01"),
  1898 => (x"41",x"43",x"47",x"4d"),
  1899 => (x"7f",x"00",x"00",x"00"),
  1900 => (x"00",x"41",x"41",x"7f"),
  1901 => (x"06",x"03",x"01",x"00"),
  1902 => (x"60",x"30",x"18",x"0c"),
  1903 => (x"41",x"00",x"00",x"40"),
  1904 => (x"00",x"7f",x"7f",x"41"),
  1905 => (x"06",x"0c",x"08",x"00"),
  1906 => (x"08",x"0c",x"06",x"03"),
  1907 => (x"80",x"80",x"80",x"00"),
  1908 => (x"80",x"80",x"80",x"80"),
  1909 => (x"00",x"00",x"00",x"00"),
  1910 => (x"00",x"04",x"07",x"03"),
  1911 => (x"74",x"20",x"00",x"00"),
  1912 => (x"78",x"7c",x"54",x"54"),
  1913 => (x"7f",x"7f",x"00",x"00"),
  1914 => (x"38",x"7c",x"44",x"44"),
  1915 => (x"7c",x"38",x"00",x"00"),
  1916 => (x"00",x"44",x"44",x"44"),
  1917 => (x"7c",x"38",x"00",x"00"),
  1918 => (x"7f",x"7f",x"44",x"44"),
  1919 => (x"7c",x"38",x"00",x"00"),
  1920 => (x"18",x"5c",x"54",x"54"),
  1921 => (x"7e",x"04",x"00",x"00"),
  1922 => (x"00",x"05",x"05",x"7f"),
  1923 => (x"bc",x"18",x"00",x"00"),
  1924 => (x"7c",x"fc",x"a4",x"a4"),
  1925 => (x"7f",x"7f",x"00",x"00"),
  1926 => (x"78",x"7c",x"04",x"04"),
  1927 => (x"00",x"00",x"00",x"00"),
  1928 => (x"00",x"40",x"7d",x"3d"),
  1929 => (x"80",x"80",x"00",x"00"),
  1930 => (x"00",x"7d",x"fd",x"80"),
  1931 => (x"7f",x"7f",x"00",x"00"),
  1932 => (x"44",x"6c",x"38",x"10"),
  1933 => (x"00",x"00",x"00",x"00"),
  1934 => (x"00",x"40",x"7f",x"3f"),
  1935 => (x"0c",x"7c",x"7c",x"00"),
  1936 => (x"78",x"7c",x"0c",x"18"),
  1937 => (x"7c",x"7c",x"00",x"00"),
  1938 => (x"78",x"7c",x"04",x"04"),
  1939 => (x"7c",x"38",x"00",x"00"),
  1940 => (x"38",x"7c",x"44",x"44"),
  1941 => (x"fc",x"fc",x"00",x"00"),
  1942 => (x"18",x"3c",x"24",x"24"),
  1943 => (x"3c",x"18",x"00",x"00"),
  1944 => (x"fc",x"fc",x"24",x"24"),
  1945 => (x"7c",x"7c",x"00",x"00"),
  1946 => (x"08",x"0c",x"04",x"04"),
  1947 => (x"5c",x"48",x"00",x"00"),
  1948 => (x"20",x"74",x"54",x"54"),
  1949 => (x"3f",x"04",x"00",x"00"),
  1950 => (x"00",x"44",x"44",x"7f"),
  1951 => (x"7c",x"3c",x"00",x"00"),
  1952 => (x"7c",x"7c",x"40",x"40"),
  1953 => (x"3c",x"1c",x"00",x"00"),
  1954 => (x"1c",x"3c",x"60",x"60"),
  1955 => (x"60",x"7c",x"3c",x"00"),
  1956 => (x"3c",x"7c",x"60",x"30"),
  1957 => (x"38",x"6c",x"44",x"00"),
  1958 => (x"44",x"6c",x"38",x"10"),
  1959 => (x"bc",x"1c",x"00",x"00"),
  1960 => (x"1c",x"3c",x"60",x"e0"),
  1961 => (x"64",x"44",x"00",x"00"),
  1962 => (x"44",x"4c",x"5c",x"74"),
  1963 => (x"08",x"08",x"00",x"00"),
  1964 => (x"41",x"41",x"77",x"3e"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"00",x"7f",x"7f"),
  1967 => (x"41",x"41",x"00",x"00"),
  1968 => (x"08",x"08",x"3e",x"77"),
  1969 => (x"01",x"01",x"02",x"00"),
  1970 => (x"01",x"02",x"02",x"03"),
  1971 => (x"7f",x"7f",x"7f",x"00"),
  1972 => (x"7f",x"7f",x"7f",x"7f"),
  1973 => (x"1c",x"08",x"08",x"00"),
  1974 => (x"7f",x"3e",x"3e",x"1c"),
  1975 => (x"3e",x"7f",x"7f",x"7f"),
  1976 => (x"08",x"1c",x"1c",x"3e"),
  1977 => (x"18",x"10",x"00",x"08"),
  1978 => (x"10",x"18",x"7c",x"7c"),
  1979 => (x"30",x"10",x"00",x"00"),
  1980 => (x"10",x"30",x"7c",x"7c"),
  1981 => (x"60",x"30",x"10",x"00"),
  1982 => (x"06",x"1e",x"78",x"60"),
  1983 => (x"3c",x"66",x"42",x"00"),
  1984 => (x"42",x"66",x"3c",x"18"),
  1985 => (x"6a",x"38",x"78",x"00"),
  1986 => (x"38",x"6c",x"c6",x"c2"),
  1987 => (x"00",x"00",x"60",x"00"),
  1988 => (x"60",x"00",x"00",x"60"),
  1989 => (x"5b",x"5e",x"0e",x"00"),
  1990 => (x"1e",x"0e",x"5d",x"5c"),
  1991 => (x"de",x"c2",x"4c",x"71"),
  1992 => (x"c0",x"4d",x"bf",x"e5"),
  1993 => (x"74",x"1e",x"c0",x"4b"),
  1994 => (x"87",x"c7",x"02",x"ab"),
  1995 => (x"c0",x"48",x"a6",x"c4"),
  1996 => (x"c4",x"87",x"c5",x"78"),
  1997 => (x"78",x"c1",x"48",x"a6"),
  1998 => (x"73",x"1e",x"66",x"c4"),
  1999 => (x"87",x"df",x"ee",x"49"),
  2000 => (x"e0",x"c0",x"86",x"c8"),
  2001 => (x"87",x"ee",x"ef",x"49"),
  2002 => (x"6a",x"4a",x"a5",x"c4"),
  2003 => (x"87",x"f0",x"f0",x"49"),
  2004 => (x"cb",x"87",x"c6",x"f1"),
  2005 => (x"c8",x"83",x"c1",x"85"),
  2006 => (x"ff",x"04",x"ab",x"b7"),
  2007 => (x"26",x"26",x"87",x"c7"),
  2008 => (x"26",x"4c",x"26",x"4d"),
  2009 => (x"1e",x"4f",x"26",x"4b"),
  2010 => (x"de",x"c2",x"4a",x"71"),
  2011 => (x"de",x"c2",x"5a",x"e9"),
  2012 => (x"78",x"c7",x"48",x"e9"),
  2013 => (x"87",x"dd",x"fe",x"49"),
  2014 => (x"73",x"1e",x"4f",x"26"),
  2015 => (x"c0",x"4a",x"71",x"1e"),
  2016 => (x"d3",x"03",x"aa",x"b7"),
  2017 => (x"c3",x"cc",x"c2",x"87"),
  2018 => (x"87",x"c4",x"05",x"bf"),
  2019 => (x"87",x"c2",x"4b",x"c1"),
  2020 => (x"cc",x"c2",x"4b",x"c0"),
  2021 => (x"87",x"c4",x"5b",x"c7"),
  2022 => (x"5a",x"c7",x"cc",x"c2"),
  2023 => (x"bf",x"c3",x"cc",x"c2"),
  2024 => (x"c1",x"9a",x"c1",x"4a"),
  2025 => (x"ec",x"49",x"a2",x"c0"),
  2026 => (x"48",x"fc",x"87",x"e8"),
  2027 => (x"bf",x"c3",x"cc",x"c2"),
  2028 => (x"87",x"ef",x"fe",x"78"),
  2029 => (x"c4",x"4a",x"71",x"1e"),
  2030 => (x"49",x"72",x"1e",x"66"),
  2031 => (x"26",x"87",x"f9",x"ea"),
  2032 => (x"ff",x"1e",x"4f",x"26"),
  2033 => (x"ff",x"c3",x"48",x"d4"),
  2034 => (x"48",x"d0",x"ff",x"78"),
  2035 => (x"ff",x"78",x"e1",x"c0"),
  2036 => (x"78",x"c1",x"48",x"d4"),
  2037 => (x"30",x"c4",x"48",x"71"),
  2038 => (x"78",x"08",x"d4",x"ff"),
  2039 => (x"c0",x"48",x"d0",x"ff"),
  2040 => (x"4f",x"26",x"78",x"e0"),
  2041 => (x"5c",x"5b",x"5e",x"0e"),
  2042 => (x"86",x"f0",x"0e",x"5d"),
  2043 => (x"c0",x"48",x"a6",x"c8"),
  2044 => (x"ec",x"4b",x"4d",x"78"),
  2045 => (x"80",x"fc",x"7e",x"bf"),
  2046 => (x"bf",x"e5",x"de",x"c2"),
  2047 => (x"4c",x"bf",x"e8",x"78"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

